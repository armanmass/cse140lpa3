-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 21 2019 00:07:27

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__22396\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu0.un165_ci_0_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un44_ci\ : std_logic;
signal \uu0.un44_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.valid_0_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_rx.idle_0_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu0.un187_ci_1\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.un143_ci_0_cascade_\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.un4_l_count_13_cascade_\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un4_l_count_16\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \CONSTANT_ONE_NET_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \resetGen.un241_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_count_2_0_4_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.un404_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.N_34\ : std_logic;
signal \uu2.N_34_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.N_31\ : std_logic;
signal \uu2.N_31_cascade_\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \INVuu2.vram_rd_clk_det_0C_net\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \G_188\ : std_logic;
signal \G_188_cascade_\ : std_logic;
signal \Lab_UT.un1_rst_0_iclkZ0\ : std_logic;
signal \G_182_cascade_\ : std_logic;
signal \G_187\ : std_logic;
signal \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\ : std_logic;
signal \G_183\ : std_logic;
signal \G_182\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu2.un28_w_addr_user_i_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_1_rep1_nesrC_net\ : std_logic;
signal \uu2.N_401\ : std_logic;
signal \uu2.N_406_cascade_\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \uu2.N_383_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\ : std_logic;
signal \uu2.bitmap_pmux_sn_i5_mux\ : std_logic;
signal \uu2.bitmap_pmux_u_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\ : std_logic;
signal \uu2.w_addr_displaying_RNI0NG56Z0Z_4\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \INVuu2.vram_rd_clk_det_1C_net\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\ : std_logic;
signal \uu2.un20_w_addr_userZ0Z_1\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \Lab_UT.dispString.N_124_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\ : std_logic;
signal \Lab_UT.didp.regrce4.LdAMtens_0\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_4\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_3\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_3\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_3\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_3\ : std_logic;
signal \Lab_UT.dispString.dOutP_1_iv_i_1_4\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\ : std_logic;
signal \G_186\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.un1_armed_2_0_iso_iZ0\ : std_logic;
signal \Lab_UT.un1_idle_4_0_iclkZ0_cascade_\ : std_logic;
signal \G_185\ : std_logic;
signal \G_185_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_117_cascade_\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\ : std_logic;
signal \G_180_cascade_\ : std_logic;
signal \G_181_cascade_\ : std_logic;
signal \G_180\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_0_cascade_\ : std_logic;
signal \Lab_UT.alarmstate_0_sqmuxa_1\ : std_logic;
signal \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\ : std_logic;
signal \G_184\ : std_logic;
signal \resetGen.escKeyZ0Z_5_cascade_\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \resetGen.escKeyZ0Z_4\ : std_logic;
signal \uu2.un28_w_addr_user_i\ : std_logic;
signal \INVuu2.w_addr_user_2C_net\ : std_logic;
signal \uu2.un51_w_data_displaying_i_a2_1\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a3_2_0\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_3C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.w_addr_displaying_RNI03P31Z0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.N_24_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.N_31_i\ : std_logic;
signal \uu2.N_26_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \Lab_UT.didp.ce_12_1\ : std_logic;
signal \Lab_UT.didp.ce_12_1_cascade_\ : std_logic;
signal \Lab_UT.didp.ce_12_3_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_1\ : std_logic;
signal \Lab_UT.dispString.N_140\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_137\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_2_2\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0_cascade_\ : std_logic;
signal \G_181\ : std_logic;
signal \G_179\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.un42_dOutP_1\ : std_logic;
signal \Lab_UT.dispString.N_95\ : std_logic;
signal \Lab_UT.didp.regrce2.LdAStens_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z8\ : std_logic;
signal \Lab_UT.dictrl.m37_N_2LZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.g1_0Z0Z_5\ : std_logic;
signal \Lab_UT.dictrl.g1_0_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_5_4_0\ : std_logic;
signal \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_5_3_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8Z0Z_3\ : std_logic;
signal \INVuu2.w_addr_displaying_ness_6C_net\ : std_logic;
signal \uu2.N_33_1\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \INVuu2.bitmap_168C_net\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux_cascade_\ : std_logic;
signal \uu2.N_14\ : std_logic;
signal \uu2.bitmap_RNI2Q8F1Z0Z_111\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.N_166\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \INVuu2.bitmap_197C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.N_149\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.N_25\ : std_logic;
signal \Lab_UT.didp.countrce1.ce_12_1_1\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.didp.countrce2.N_93\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\ : std_logic;
signal \Lab_UT.didp.countrce2.N_96_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.un24_ce_3\ : std_logic;
signal \Lab_UT.dispString.N_143\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_0\ : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2\ : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\ : std_logic;
signal \Lab_UT.didp.N_90\ : std_logic;
signal \Lab_UT.LdSones_i_4\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.state_ret_8_ess\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1\ : std_logic;
signal \Lab_UT.didp.regrce1.LdASones_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_a5_1_0_cascade_\ : std_logic;
signal \Lab_UT.i8_mux_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_sn\ : std_logic;
signal \Lab_UT.dictrl.g1_1_0_1_cascade_\ : std_logic;
signal \Lab_UT.g1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_rn_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_1\ : std_logic;
signal \Lab_UT.dictrl.g2Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g0_6_3_0\ : std_logic;
signal \Lab_UT.dictrl.m13_out_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_18_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_5\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_4\ : std_logic;
signal \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_11\ : std_logic;
signal \Lab_UT.dictrl.m34Z0Z_1_cascade_\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal \Lab_UT.dictrl.m22Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux_1\ : std_logic;
signal \Lab_UT.dictrl.g1_1_0_0\ : std_logic;
signal \Lab_UT.dictrl.m22Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g1_1_0\ : std_logic;
signal \Lab_UT.dictrl.g1_rn_0\ : std_logic;
signal \Lab_UT.dictrl.m34Z0Z_1\ : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal \Lab_UT.dictrl.g1_1_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_1Z0Z_5\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \uu2.N_40\ : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_8C_net\ : std_logic;
signal \uu2.N_37\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.N_45\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_36\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmap_pmux_20_ns_1\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.bitmap_pmux_26_bm_1\ : std_logic;
signal \uu2.bitmap_RNIP2JO1Z0Z_34\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.min1_0\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.min1_3\ : std_logic;
signal \Lab_UT.sec1_3\ : std_logic;
signal \Lab_UT.sec1_0\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \uu2.bitmap_pmux_17_ns_1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.bitmap_pmux_16_ns_1\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \Lab_UT.min2_0\ : std_logic;
signal \Lab_UT.min2_3\ : std_logic;
signal \Lab_UT.min2_2\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \INVuu2.bitmap_215C_net\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.sec1_1\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.min1_1\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.sec1_2\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal \Lab_UT.didp.countrce1.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0\ : std_logic;
signal \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\ : std_logic;
signal \Lab_UT.min2_1\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.min1_2\ : std_logic;
signal \Lab_UT.didp.regrce3.LdAMones_0\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.dispString.N_118_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_1\ : std_logic;
signal \Lab_UT.dispString.N_145\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMones_1\ : std_logic;
signal \Lab_UT.LdAMones\ : std_logic;
signal \Lab_UT.LdAMones_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_rn_0\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_57_1\ : std_logic;
signal \Lab_UT.dictrl.N_55_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_sn\ : std_logic;
signal \Lab_UT.dictrl.un15_loadalarm_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.loadalarm_0_0\ : std_logic;
signal \Lab_UT.LdAStens\ : std_logic;
signal \Lab_UT.dictrl.N_22\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_1\ : std_logic;
signal \Lab_UT.dictrl.g2_0_0\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_2\ : std_logic;
signal \Lab_UT.dictrl.N_20_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_22_0_0\ : std_logic;
signal \Lab_UT.next_state_0\ : std_logic;
signal \Lab_UT.next_state_1_0_0_1_cascade_\ : std_logic;
signal \Lab_UT.next_state_2\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.didp.g0_0_2Z0Z_1\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.didp.g0_0Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state6\ : std_logic;
signal \Lab_UT.dictrl.N_20_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m34_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_26_0\ : std_logic;
signal \Lab_UT.dictrl.m34_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_60_0_0\ : std_logic;
signal \Lab_UT.dictrl.m19_1\ : std_logic;
signal \N_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_59_1_0\ : std_logic;
signal \Lab_UT.dictrl.i8_mux_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13\ : std_logic;
signal \Lab_UT.dictrl.m22_xZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m22Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_18\ : std_logic;
signal m7_a0 : std_logic;
signal \Lab_UT.dictrl.state_fast_0\ : std_logic;
signal \buart__rx_shifter_fast_4\ : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_6_3\ : std_logic;
signal \Lab_UT.dictrl.gZ0Z2\ : std_logic;
signal \Lab_UT.dictrl.g0_6_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_1\ : std_logic;
signal \Lab_UT.dictrl.N_57_0\ : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal \Lab_UT.dictrl.g1_0_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0_xZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.g0_5Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.g0_5_3\ : std_logic;
signal \Lab_UT.dictrl.g1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_55_0\ : std_logic;
signal \Lab_UT.dictrl.g0_3_4_cascade_\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal \Lab_UT.dictrl.N_72_mux_0\ : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \Lab_UT.dictrl.g0_3_3\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.un3_w_addr_user_4_cascade_\ : std_logic;
signal \uu2.un3_w_addr_user_5\ : std_logic;
signal \uu2.un3_w_addr_user\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.un404_ci_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.un426_ci_3\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.vbuf_w_addr_user.un448_ci_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.w_addr_user_RNI43E87Z0Z_4\ : std_logic;
signal \uu2.N_44\ : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_8\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \INVuu2.w_addr_displaying_7C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmap_pmux_19_ns_1\ : std_logic;
signal \Lab_UT.sec2_0\ : std_logic;
signal \Lab_UT.sec2_3\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.N_152_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \uu2.bitmap_RNIM5E21Z0Z_314\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.reset_12_1_3\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_144\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.sec2_2\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMtens_0\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.loadalarm_0\ : std_logic;
signal \Lab_UT.sec2_1\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.countrce4.un13_qPone\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2\ : std_logic;
signal \uu0_sec_clkD\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \oneSecStrb_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_102\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.dictrl.state_i_3_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_2_fast\ : std_logic;
signal \Lab_UT.dictrl.N_20\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_1\ : std_logic;
signal \Lab_UT.dictrl.m19_1_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_3\ : std_logic;
signal \Lab_UT.next_state_1\ : std_logic;
signal \Lab_UT.dictrl.next_state66_2\ : std_logic;
signal \Lab_UT.bu_rx_data_rdy_0\ : std_logic;
signal \Lab_UT.state_i_4_3\ : std_logic;
signal \Lab_UT.dictrl.dicRun_1\ : std_logic;
signal \Lab_UT.state_2\ : std_logic;
signal \Lab_UT.LdASones\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.g1_4_0\ : std_logic;
signal \Lab_UT.dictrl.g1_5_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_4_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_0\ : std_logic;
signal \shifter_1_rep1_RNI0FPF_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_33_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_1\ : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_1\ : std_logic;
signal \N_15_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_20_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.g0_0\ : std_logic;
signal \Lab_UT.dictrl.N_15_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_60_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0\ : std_logic;
signal \Lab_UT.un1_next_state66_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_60\ : std_logic;
signal \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\ : std_logic;
signal \Lab_UT.dicLdSones_1\ : std_logic;
signal \G_6_0_a6_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_0_1\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_1_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m13_out\ : std_logic;
signal \Lab_UT.dictrl.N_15_0\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux\ : std_logic;
signal \Lab_UT.dictrl.N_59\ : std_logic;
signal \Lab_UT.dictrl.N_8_0\ : std_logic;
signal \Lab_UT.dictrl.i8_mux\ : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal \Lab_UT.dictrl.state_0_rep1\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_3\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_5Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.i9_mux\ : std_logic;
signal \Lab_UT_dictrl_state_1\ : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal \Lab_UT.dictrl.N_67_mux\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_3\ : std_logic;
signal \G_6_0_a6_3_3_cascade_\ : std_logic;
signal \Lab_UT.stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_12\ : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal \N_63_mux\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_3_rep2 : std_logic;
signal \N_14_0\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_2 : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal rst_g : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal clk_g : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__9780\&\N__10050\&\N__10029\&\N__10482\&\N__10116\&\N__9759\&\N__10275\&\N__10248\&\N__10215\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__10533\&\N__11826\&\N__11865\&\N__11838\&\N__11850\&\N__16056\&\N__21627\&\N__20241\&\N__9582\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__9999\&'0'&\N__9993\&'0'&\N__9966\&'0'&\N__9978\&'0'&\N__21855\&'0'&\N__9972\&'0'&\N__10281\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__8085\,
            RESETB => \N__11095\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22269\,
            RE => \N__11100\,
            WCLKE => \N__10517\,
            WCLK => \N__22268\,
            WE => \N__10521\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22396\,
            DIN => \N__22395\,
            DOUT => \N__22394\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22396\,
            PADOUT => \N__22395\,
            PADIN => \N__22394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22387\,
            DIN => \N__22386\,
            DOUT => \N__22385\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22387\,
            PADOUT => \N__22386\,
            PADIN => \N__22385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22378\,
            DIN => \N__22377\,
            DOUT => \N__22376\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22378\,
            PADOUT => \N__22377\,
            PADIN => \N__22376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22369\,
            DIN => \N__22368\,
            DOUT => \N__22367\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__22369\,
            PADOUT => \N__22368\,
            PADIN => \N__22367\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__22223\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22360\,
            DIN => \N__22359\,
            DOUT => \N__22358\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22360\,
            PADOUT => \N__22359\,
            PADIN => \N__22358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22351\,
            DIN => \N__22350\,
            DOUT => \N__22349\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22351\,
            PADOUT => \N__22350\,
            PADIN => \N__22349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22342\,
            DIN => \N__22341\,
            DOUT => \N__22340\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22342\,
            PADOUT => \N__22341\,
            PADIN => \N__22340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22333\,
            DIN => \N__22332\,
            DOUT => \N__22331\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22333\,
            PADOUT => \N__22332\,
            PADIN => \N__22331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22324\,
            DIN => \N__22323\,
            DOUT => \N__22322\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22324\,
            PADOUT => \N__22323\,
            PADIN => \N__22322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22315\,
            DIN => \N__22314\,
            DOUT => \N__22313\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22315\,
            PADOUT => \N__22314\,
            PADIN => \N__22313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5423\ : InMux
    port map (
            O => \N__22296\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__5422\ : InMux
    port map (
            O => \N__22293\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__5421\ : InMux
    port map (
            O => \N__22290\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__5420\ : InMux
    port map (
            O => \N__22287\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__5419\ : InMux
    port map (
            O => \N__22284\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__22281\,
            I => \N__22278\
        );

    \I__5417\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22275\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__22275\,
            I => \N__22185\
        );

    \I__5415\ : ClkMux
    port map (
            O => \N__22274\,
            I => \N__22008\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__22273\,
            I => \N__22008\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__22272\,
            I => \N__22008\
        );

    \I__5412\ : ClkMux
    port map (
            O => \N__22271\,
            I => \N__22008\
        );

    \I__5411\ : ClkMux
    port map (
            O => \N__22270\,
            I => \N__22008\
        );

    \I__5410\ : ClkMux
    port map (
            O => \N__22269\,
            I => \N__22008\
        );

    \I__5409\ : ClkMux
    port map (
            O => \N__22268\,
            I => \N__22008\
        );

    \I__5408\ : ClkMux
    port map (
            O => \N__22267\,
            I => \N__22008\
        );

    \I__5407\ : ClkMux
    port map (
            O => \N__22266\,
            I => \N__22008\
        );

    \I__5406\ : ClkMux
    port map (
            O => \N__22265\,
            I => \N__22008\
        );

    \I__5405\ : ClkMux
    port map (
            O => \N__22264\,
            I => \N__22008\
        );

    \I__5404\ : ClkMux
    port map (
            O => \N__22263\,
            I => \N__22008\
        );

    \I__5403\ : ClkMux
    port map (
            O => \N__22262\,
            I => \N__22008\
        );

    \I__5402\ : ClkMux
    port map (
            O => \N__22261\,
            I => \N__22008\
        );

    \I__5401\ : ClkMux
    port map (
            O => \N__22260\,
            I => \N__22008\
        );

    \I__5400\ : ClkMux
    port map (
            O => \N__22259\,
            I => \N__22008\
        );

    \I__5399\ : ClkMux
    port map (
            O => \N__22258\,
            I => \N__22008\
        );

    \I__5398\ : ClkMux
    port map (
            O => \N__22257\,
            I => \N__22008\
        );

    \I__5397\ : ClkMux
    port map (
            O => \N__22256\,
            I => \N__22008\
        );

    \I__5396\ : ClkMux
    port map (
            O => \N__22255\,
            I => \N__22008\
        );

    \I__5395\ : ClkMux
    port map (
            O => \N__22254\,
            I => \N__22008\
        );

    \I__5394\ : ClkMux
    port map (
            O => \N__22253\,
            I => \N__22008\
        );

    \I__5393\ : ClkMux
    port map (
            O => \N__22252\,
            I => \N__22008\
        );

    \I__5392\ : ClkMux
    port map (
            O => \N__22251\,
            I => \N__22008\
        );

    \I__5391\ : ClkMux
    port map (
            O => \N__22250\,
            I => \N__22008\
        );

    \I__5390\ : ClkMux
    port map (
            O => \N__22249\,
            I => \N__22008\
        );

    \I__5389\ : ClkMux
    port map (
            O => \N__22248\,
            I => \N__22008\
        );

    \I__5388\ : ClkMux
    port map (
            O => \N__22247\,
            I => \N__22008\
        );

    \I__5387\ : ClkMux
    port map (
            O => \N__22246\,
            I => \N__22008\
        );

    \I__5386\ : ClkMux
    port map (
            O => \N__22245\,
            I => \N__22008\
        );

    \I__5385\ : ClkMux
    port map (
            O => \N__22244\,
            I => \N__22008\
        );

    \I__5384\ : ClkMux
    port map (
            O => \N__22243\,
            I => \N__22008\
        );

    \I__5383\ : ClkMux
    port map (
            O => \N__22242\,
            I => \N__22008\
        );

    \I__5382\ : ClkMux
    port map (
            O => \N__22241\,
            I => \N__22008\
        );

    \I__5381\ : ClkMux
    port map (
            O => \N__22240\,
            I => \N__22008\
        );

    \I__5380\ : ClkMux
    port map (
            O => \N__22239\,
            I => \N__22008\
        );

    \I__5379\ : ClkMux
    port map (
            O => \N__22238\,
            I => \N__22008\
        );

    \I__5378\ : ClkMux
    port map (
            O => \N__22237\,
            I => \N__22008\
        );

    \I__5377\ : ClkMux
    port map (
            O => \N__22236\,
            I => \N__22008\
        );

    \I__5376\ : ClkMux
    port map (
            O => \N__22235\,
            I => \N__22008\
        );

    \I__5375\ : ClkMux
    port map (
            O => \N__22234\,
            I => \N__22008\
        );

    \I__5374\ : ClkMux
    port map (
            O => \N__22233\,
            I => \N__22008\
        );

    \I__5373\ : ClkMux
    port map (
            O => \N__22232\,
            I => \N__22008\
        );

    \I__5372\ : ClkMux
    port map (
            O => \N__22231\,
            I => \N__22008\
        );

    \I__5371\ : ClkMux
    port map (
            O => \N__22230\,
            I => \N__22008\
        );

    \I__5370\ : ClkMux
    port map (
            O => \N__22229\,
            I => \N__22008\
        );

    \I__5369\ : ClkMux
    port map (
            O => \N__22228\,
            I => \N__22008\
        );

    \I__5368\ : ClkMux
    port map (
            O => \N__22227\,
            I => \N__22008\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22226\,
            I => \N__22008\
        );

    \I__5366\ : ClkMux
    port map (
            O => \N__22225\,
            I => \N__22008\
        );

    \I__5365\ : ClkMux
    port map (
            O => \N__22224\,
            I => \N__22008\
        );

    \I__5364\ : ClkMux
    port map (
            O => \N__22223\,
            I => \N__22008\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22222\,
            I => \N__22008\
        );

    \I__5362\ : ClkMux
    port map (
            O => \N__22221\,
            I => \N__22008\
        );

    \I__5361\ : ClkMux
    port map (
            O => \N__22220\,
            I => \N__22008\
        );

    \I__5360\ : ClkMux
    port map (
            O => \N__22219\,
            I => \N__22008\
        );

    \I__5359\ : ClkMux
    port map (
            O => \N__22218\,
            I => \N__22008\
        );

    \I__5358\ : ClkMux
    port map (
            O => \N__22217\,
            I => \N__22008\
        );

    \I__5357\ : ClkMux
    port map (
            O => \N__22216\,
            I => \N__22008\
        );

    \I__5356\ : ClkMux
    port map (
            O => \N__22215\,
            I => \N__22008\
        );

    \I__5355\ : ClkMux
    port map (
            O => \N__22214\,
            I => \N__22008\
        );

    \I__5354\ : ClkMux
    port map (
            O => \N__22213\,
            I => \N__22008\
        );

    \I__5353\ : ClkMux
    port map (
            O => \N__22212\,
            I => \N__22008\
        );

    \I__5352\ : ClkMux
    port map (
            O => \N__22211\,
            I => \N__22008\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__22210\,
            I => \N__22008\
        );

    \I__5350\ : ClkMux
    port map (
            O => \N__22209\,
            I => \N__22008\
        );

    \I__5349\ : ClkMux
    port map (
            O => \N__22208\,
            I => \N__22008\
        );

    \I__5348\ : ClkMux
    port map (
            O => \N__22207\,
            I => \N__22008\
        );

    \I__5347\ : ClkMux
    port map (
            O => \N__22206\,
            I => \N__22008\
        );

    \I__5346\ : ClkMux
    port map (
            O => \N__22205\,
            I => \N__22008\
        );

    \I__5345\ : ClkMux
    port map (
            O => \N__22204\,
            I => \N__22008\
        );

    \I__5344\ : ClkMux
    port map (
            O => \N__22203\,
            I => \N__22008\
        );

    \I__5343\ : ClkMux
    port map (
            O => \N__22202\,
            I => \N__22008\
        );

    \I__5342\ : ClkMux
    port map (
            O => \N__22201\,
            I => \N__22008\
        );

    \I__5341\ : ClkMux
    port map (
            O => \N__22200\,
            I => \N__22008\
        );

    \I__5340\ : ClkMux
    port map (
            O => \N__22199\,
            I => \N__22008\
        );

    \I__5339\ : ClkMux
    port map (
            O => \N__22198\,
            I => \N__22008\
        );

    \I__5338\ : ClkMux
    port map (
            O => \N__22197\,
            I => \N__22008\
        );

    \I__5337\ : ClkMux
    port map (
            O => \N__22196\,
            I => \N__22008\
        );

    \I__5336\ : ClkMux
    port map (
            O => \N__22195\,
            I => \N__22008\
        );

    \I__5335\ : ClkMux
    port map (
            O => \N__22194\,
            I => \N__22008\
        );

    \I__5334\ : ClkMux
    port map (
            O => \N__22193\,
            I => \N__22008\
        );

    \I__5333\ : ClkMux
    port map (
            O => \N__22192\,
            I => \N__22008\
        );

    \I__5332\ : ClkMux
    port map (
            O => \N__22191\,
            I => \N__22008\
        );

    \I__5331\ : ClkMux
    port map (
            O => \N__22190\,
            I => \N__22008\
        );

    \I__5330\ : ClkMux
    port map (
            O => \N__22189\,
            I => \N__22008\
        );

    \I__5329\ : ClkMux
    port map (
            O => \N__22188\,
            I => \N__22008\
        );

    \I__5328\ : Glb2LocalMux
    port map (
            O => \N__22185\,
            I => \N__22008\
        );

    \I__5327\ : GlobalMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__5326\ : gio2CtrlBuf
    port map (
            O => \N__22005\,
            I => clk_g
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__22002\,
            I => \N__21999\
        );

    \I__5324\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21993\
        );

    \I__5323\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21993\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__21993\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__5320\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21981\
        );

    \I__5319\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21981\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__21981\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__21978\,
            I => \N__21974\
        );

    \I__5316\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21971\
        );

    \I__5315\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21968\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__21971\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__21968\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__5312\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21957\
        );

    \I__5311\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21957\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__21957\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__5309\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21949\
        );

    \I__5308\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21944\
        );

    \I__5307\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21944\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__21949\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__21944\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__21939\,
            I => \N__21934\
        );

    \I__5303\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21928\
        );

    \I__5302\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21928\
        );

    \I__5301\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21923\
        );

    \I__5300\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21923\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__21928\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__21923\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__21918\,
            I => \N__21914\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__21917\,
            I => \N__21911\
        );

    \I__5295\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21906\
        );

    \I__5294\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21906\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__21906\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__5292\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__21900\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__5290\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21887\
        );

    \I__5289\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21887\
        );

    \I__5288\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21887\
        );

    \I__5287\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21884\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__21887\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__21884\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__5284\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__5282\ : Span4Mux_s3_v
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__21870\,
            I => \N__21865\
        );

    \I__5280\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21860\
        );

    \I__5279\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21860\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__21865\,
            I => \L3_tx_data_2\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__21860\,
            I => \L3_tx_data_2\
        );

    \I__5276\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__5274\ : Span4Mux_s0_v
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__21843\,
            I => \uu2.mem0.w_data_2\
        );

    \I__5271\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21833\
        );

    \I__5270\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21830\
        );

    \I__5269\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21825\
        );

    \I__5268\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21825\
        );

    \I__5267\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21822\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21819\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21814\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21814\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__21822\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5262\ : Odrv12
    port map (
            O => \N__21819\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__21814\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5260\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21796\
        );

    \I__5259\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21796\
        );

    \I__5258\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21796\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__21804\,
            I => \N__21793\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__21803\,
            I => \N__21790\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21782\
        );

    \I__5254\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21773\
        );

    \I__5253\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21773\
        );

    \I__5252\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21773\
        );

    \I__5251\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21773\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__21787\,
            I => \N__21769\
        );

    \I__5249\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21761\
        );

    \I__5248\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21758\
        );

    \I__5247\ : Span4Mux_s2_v
    port map (
            O => \N__21782\,
            I => \N__21755\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21752\
        );

    \I__5245\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21749\
        );

    \I__5244\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21735\
        );

    \I__5243\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21735\
        );

    \I__5242\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21735\
        );

    \I__5241\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21735\
        );

    \I__5240\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21735\
        );

    \I__5239\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21735\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21730\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21730\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__21755\,
            I => \N__21725\
        );

    \I__5235\ : Span4Mux_s2_v
    port map (
            O => \N__21752\,
            I => \N__21725\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21722\
        );

    \I__5233\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21719\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21716\
        );

    \I__5231\ : Span4Mux_s2_v
    port map (
            O => \N__21730\,
            I => \N__21713\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__21725\,
            I => \N__21708\
        );

    \I__5229\ : Span4Mux_v
    port map (
            O => \N__21722\,
            I => \N__21708\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21705\
        );

    \I__5227\ : Span4Mux_s2_v
    port map (
            O => \N__21716\,
            I => \N__21700\
        );

    \I__5226\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21700\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__21708\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5224\ : Odrv12
    port map (
            O => \N__21705\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__21700\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21689\
        );

    \I__5221\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21685\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21682\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__21688\,
            I => \N__21679\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__21685\,
            I => \N__21667\
        );

    \I__5217\ : Span4Mux_s2_v
    port map (
            O => \N__21682\,
            I => \N__21664\
        );

    \I__5216\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21655\
        );

    \I__5215\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21655\
        );

    \I__5214\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21655\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21655\
        );

    \I__5212\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21650\
        );

    \I__5211\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21650\
        );

    \I__5210\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21641\
        );

    \I__5209\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21641\
        );

    \I__5208\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21641\
        );

    \I__5207\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21641\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__21667\,
            I => \N__21638\
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__21664\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__21655\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__21650\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__21641\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__21638\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__5199\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21618\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__5196\ : Span4Mux_h
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__21612\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__5194\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21606\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__21606\,
            I => \buart.Z_tx.un1_bitcount_c2\
        );

    \I__5192\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21599\
        );

    \I__5191\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__21599\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__21596\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__21591\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__21588\,
            I => \N__21585\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21577\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21574\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21565\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21565\
        );

    \I__5182\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21565\
        );

    \I__5181\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21565\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21577\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21574\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__21565\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__5177\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21552\
        );

    \I__5176\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21545\
        );

    \I__5175\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21545\
        );

    \I__5174\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21545\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__21552\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__21545\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21535\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21530\
        );

    \I__5169\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21530\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21535\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__21530\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__5165\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21513\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21513\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21506\
        );

    \I__5162\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21506\
        );

    \I__5161\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21506\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__21513\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21506\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21498\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__21498\,
            I => \buart.Z_tx.un1_bitcount_c3\
        );

    \I__5156\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21487\
        );

    \I__5155\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21487\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__21493\,
            I => \N__21483\
        );

    \I__5153\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21477\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__21487\,
            I => \N__21474\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21469\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21469\
        );

    \I__5149\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21462\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21459\
        );

    \I__5147\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21456\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__21477\,
            I => \N__21449\
        );

    \I__5145\ : Span4Mux_h
    port map (
            O => \N__21474\,
            I => \N__21449\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__21469\,
            I => \N__21449\
        );

    \I__5143\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21446\
        );

    \I__5142\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21439\
        );

    \I__5141\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21439\
        );

    \I__5140\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21439\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21432\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21429\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21424\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__21449\,
            I => \N__21424\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21446\,
            I => \N__21419\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21439\,
            I => \N__21419\
        );

    \I__5133\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21410\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21410\
        );

    \I__5131\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21410\
        );

    \I__5130\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21410\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__21432\,
            I => \N__21407\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__21429\,
            I => \N_63_mux\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__21424\,
            I => \N_63_mux\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__21419\,
            I => \N_63_mux\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N_63_mux\
        );

    \I__5124\ : Odrv4
    port map (
            O => \N__21407\,
            I => \N_63_mux\
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__21396\,
            I => \N__21392\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21386\
        );

    \I__5121\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21383\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__21391\,
            I => \N__21380\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21374\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21371\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__21386\,
            I => \N__21368\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21365\
        );

    \I__5115\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21362\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__21379\,
            I => \N__21359\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21356\
        );

    \I__5112\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21353\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21349\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21340\
        );

    \I__5109\ : Span4Mux_s3_h
    port map (
            O => \N__21368\,
            I => \N__21340\
        );

    \I__5108\ : Span4Mux_s3_h
    port map (
            O => \N__21365\,
            I => \N__21340\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21340\
        );

    \I__5106\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21337\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21330\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21330\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21327\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__21349\,
            I => \N__21322\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__21340\,
            I => \N__21322\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21319\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21316\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21309\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__21330\,
            I => \N__21303\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__21327\,
            I => \N__21300\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__21322\,
            I => \N__21297\
        );

    \I__5094\ : Span4Mux_v
    port map (
            O => \N__21319\,
            I => \N__21292\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21292\
        );

    \I__5092\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21287\
        );

    \I__5091\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21287\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21282\
        );

    \I__5089\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21282\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21279\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21274\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21274\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21271\
        );

    \I__5084\ : Span4Mux_v
    port map (
            O => \N__21303\,
            I => \N__21268\
        );

    \I__5083\ : Span4Mux_h
    port map (
            O => \N__21300\,
            I => \N__21263\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__21297\,
            I => \N__21263\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__21292\,
            I => \N__21258\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21258\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21282\,
            I => \N__21255\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21279\,
            I => \N__21252\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21274\,
            I => bu_rx_data_1
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__21271\,
            I => bu_rx_data_1
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__21268\,
            I => bu_rx_data_1
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__21263\,
            I => bu_rx_data_1
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__21258\,
            I => bu_rx_data_1
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__21255\,
            I => bu_rx_data_1
        );

    \I__5071\ : Odrv12
    port map (
            O => \N__21252\,
            I => bu_rx_data_1
        );

    \I__5070\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21224\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21224\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21218\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21218\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21215\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21207\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21207\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21202\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21202\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21199\
        );

    \I__5060\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21196\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21193\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21190\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21187\
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__21213\,
            I => \N__21184\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21181\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21176\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21176\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__21199\,
            I => \N__21165\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21165\
        );

    \I__5050\ : Span4Mux_s3_h
    port map (
            O => \N__21193\,
            I => \N__21165\
        );

    \I__5049\ : Span4Mux_s3_v
    port map (
            O => \N__21190\,
            I => \N__21165\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21165\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21162\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__21181\,
            I => bu_rx_data_3_rep2
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__21176\,
            I => bu_rx_data_3_rep2
        );

    \I__5044\ : Odrv4
    port map (
            O => \N__21165\,
            I => bu_rx_data_3_rep2
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21162\,
            I => bu_rx_data_3_rep2
        );

    \I__5042\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21147\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21147\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__5039\ : Odrv12
    port map (
            O => \N__21144\,
            I => \N_14_0\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21137\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21131\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21137\,
            I => \N__21128\
        );

    \I__5035\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21125\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \N__21122\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21118\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21131\,
            I => \N__21108\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__21128\,
            I => \N__21108\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21108\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21105\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21101\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21118\,
            I => \N__21098\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21088\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21085\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21081\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__21108\,
            I => \N__21078\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21105\,
            I => \N__21075\
        );

    \I__5021\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21072\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21069\
        );

    \I__5019\ : Span4Mux_v
    port map (
            O => \N__21098\,
            I => \N__21066\
        );

    \I__5018\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21061\
        );

    \I__5017\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21061\
        );

    \I__5016\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21058\
        );

    \I__5015\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21055\
        );

    \I__5014\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21051\
        );

    \I__5013\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21048\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21045\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21039\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21039\
        );

    \I__5009\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21036\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__21081\,
            I => \N__21033\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__21078\,
            I => \N__21030\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__21075\,
            I => \N__21025\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21025\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__21069\,
            I => \N__21022\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__21066\,
            I => \N__21015\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21015\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21015\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21012\
        );

    \I__4999\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21009\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21004\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21004\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__21045\,
            I => \N__21001\
        );

    \I__4995\ : InMux
    port map (
            O => \N__21044\,
            I => \N__20998\
        );

    \I__4994\ : Span12Mux_v
    port map (
            O => \N__21039\,
            I => \N__20995\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21036\,
            I => \N__20988\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__21033\,
            I => \N__20988\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__21030\,
            I => \N__20988\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__21025\,
            I => \N__20985\
        );

    \I__4989\ : Span4Mux_v
    port map (
            O => \N__21022\,
            I => \N__20980\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__21015\,
            I => \N__20980\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__21012\,
            I => \N__20971\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__20971\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__21004\,
            I => \N__20971\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20971\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__20998\,
            I => bu_rx_data_3
        );

    \I__4982\ : Odrv12
    port map (
            O => \N__20995\,
            I => bu_rx_data_3
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__20988\,
            I => bu_rx_data_3
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__20985\,
            I => bu_rx_data_3
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__20980\,
            I => bu_rx_data_3
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__20971\,
            I => bu_rx_data_3
        );

    \I__4977\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20953\
        );

    \I__4976\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20950\
        );

    \I__4975\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20947\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20940\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__20950\,
            I => \N__20940\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__20947\,
            I => \N__20937\
        );

    \I__4971\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20934\
        );

    \I__4970\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20929\
        );

    \I__4969\ : Span4Mux_v
    port map (
            O => \N__20940\,
            I => \N__20919\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__20937\,
            I => \N__20919\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20919\
        );

    \I__4966\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20916\
        );

    \I__4965\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20913\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__20929\,
            I => \N__20910\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__20928\,
            I => \N__20905\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__20927\,
            I => \N__20901\
        );

    \I__4961\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20897\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__20919\,
            I => \N__20894\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20889\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__20913\,
            I => \N__20889\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__20910\,
            I => \N__20886\
        );

    \I__4956\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20883\
        );

    \I__4955\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20880\
        );

    \I__4954\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20875\
        );

    \I__4953\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20875\
        );

    \I__4952\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20871\
        );

    \I__4951\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20868\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__20897\,
            I => \N__20865\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__20894\,
            I => \N__20862\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__20889\,
            I => \N__20858\
        );

    \I__4947\ : Span4Mux_v
    port map (
            O => \N__20886\,
            I => \N__20849\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20849\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20849\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__20875\,
            I => \N__20849\
        );

    \I__4943\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20843\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20840\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__20868\,
            I => \N__20837\
        );

    \I__4940\ : Span12Mux_s8_v
    port map (
            O => \N__20865\,
            I => \N__20834\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__20862\,
            I => \N__20831\
        );

    \I__4938\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20828\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__20858\,
            I => \N__20823\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__20849\,
            I => \N__20823\
        );

    \I__4935\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20816\
        );

    \I__4934\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20816\
        );

    \I__4933\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20816\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20843\,
            I => \N__20811\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__20840\,
            I => \N__20811\
        );

    \I__4930\ : Odrv12
    port map (
            O => \N__20837\,
            I => bu_rx_data_2
        );

    \I__4929\ : Odrv12
    port map (
            O => \N__20834\,
            I => bu_rx_data_2
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__20831\,
            I => bu_rx_data_2
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__20828\,
            I => bu_rx_data_2
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__20823\,
            I => bu_rx_data_2
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__20816\,
            I => bu_rx_data_2
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__20811\,
            I => bu_rx_data_2
        );

    \I__4923\ : CEMux
    port map (
            O => \N__20796\,
            I => \N__20772\
        );

    \I__4922\ : CEMux
    port map (
            O => \N__20795\,
            I => \N__20772\
        );

    \I__4921\ : CEMux
    port map (
            O => \N__20794\,
            I => \N__20772\
        );

    \I__4920\ : CEMux
    port map (
            O => \N__20793\,
            I => \N__20772\
        );

    \I__4919\ : CEMux
    port map (
            O => \N__20792\,
            I => \N__20772\
        );

    \I__4918\ : CEMux
    port map (
            O => \N__20791\,
            I => \N__20772\
        );

    \I__4917\ : CEMux
    port map (
            O => \N__20790\,
            I => \N__20772\
        );

    \I__4916\ : CEMux
    port map (
            O => \N__20789\,
            I => \N__20772\
        );

    \I__4915\ : GlobalMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__4914\ : gio2CtrlBuf
    port map (
            O => \N__20769\,
            I => \buart.Z_rx.sample_g\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__20766\,
            I => \N__20758\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__20765\,
            I => \N__20751\
        );

    \I__4911\ : InMux
    port map (
            O => \N__20764\,
            I => \N__20743\
        );

    \I__4910\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20740\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20737\
        );

    \I__4908\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20734\
        );

    \I__4907\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20731\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20728\
        );

    \I__4905\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20723\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20723\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20720\
        );

    \I__4902\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20717\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20714\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20711\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20708\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20703\
        );

    \I__4897\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20703\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20743\,
            I => \N__20700\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20655\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20652\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__20734\,
            I => \N__20649\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20646\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__20728\,
            I => \N__20643\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__20723\,
            I => \N__20640\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__20720\,
            I => \N__20637\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__20717\,
            I => \N__20634\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__20714\,
            I => \N__20631\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20614\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20708\,
            I => \N__20611\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__20703\,
            I => \N__20608\
        );

    \I__4883\ : Glb2LocalMux
    port map (
            O => \N__20700\,
            I => \N__20469\
        );

    \I__4882\ : SRMux
    port map (
            O => \N__20699\,
            I => \N__20469\
        );

    \I__4881\ : SRMux
    port map (
            O => \N__20698\,
            I => \N__20469\
        );

    \I__4880\ : SRMux
    port map (
            O => \N__20697\,
            I => \N__20469\
        );

    \I__4879\ : SRMux
    port map (
            O => \N__20696\,
            I => \N__20469\
        );

    \I__4878\ : SRMux
    port map (
            O => \N__20695\,
            I => \N__20469\
        );

    \I__4877\ : SRMux
    port map (
            O => \N__20694\,
            I => \N__20469\
        );

    \I__4876\ : SRMux
    port map (
            O => \N__20693\,
            I => \N__20469\
        );

    \I__4875\ : SRMux
    port map (
            O => \N__20692\,
            I => \N__20469\
        );

    \I__4874\ : SRMux
    port map (
            O => \N__20691\,
            I => \N__20469\
        );

    \I__4873\ : SRMux
    port map (
            O => \N__20690\,
            I => \N__20469\
        );

    \I__4872\ : SRMux
    port map (
            O => \N__20689\,
            I => \N__20469\
        );

    \I__4871\ : SRMux
    port map (
            O => \N__20688\,
            I => \N__20469\
        );

    \I__4870\ : SRMux
    port map (
            O => \N__20687\,
            I => \N__20469\
        );

    \I__4869\ : SRMux
    port map (
            O => \N__20686\,
            I => \N__20469\
        );

    \I__4868\ : SRMux
    port map (
            O => \N__20685\,
            I => \N__20469\
        );

    \I__4867\ : SRMux
    port map (
            O => \N__20684\,
            I => \N__20469\
        );

    \I__4866\ : SRMux
    port map (
            O => \N__20683\,
            I => \N__20469\
        );

    \I__4865\ : SRMux
    port map (
            O => \N__20682\,
            I => \N__20469\
        );

    \I__4864\ : SRMux
    port map (
            O => \N__20681\,
            I => \N__20469\
        );

    \I__4863\ : SRMux
    port map (
            O => \N__20680\,
            I => \N__20469\
        );

    \I__4862\ : SRMux
    port map (
            O => \N__20679\,
            I => \N__20469\
        );

    \I__4861\ : SRMux
    port map (
            O => \N__20678\,
            I => \N__20469\
        );

    \I__4860\ : SRMux
    port map (
            O => \N__20677\,
            I => \N__20469\
        );

    \I__4859\ : SRMux
    port map (
            O => \N__20676\,
            I => \N__20469\
        );

    \I__4858\ : SRMux
    port map (
            O => \N__20675\,
            I => \N__20469\
        );

    \I__4857\ : SRMux
    port map (
            O => \N__20674\,
            I => \N__20469\
        );

    \I__4856\ : SRMux
    port map (
            O => \N__20673\,
            I => \N__20469\
        );

    \I__4855\ : SRMux
    port map (
            O => \N__20672\,
            I => \N__20469\
        );

    \I__4854\ : SRMux
    port map (
            O => \N__20671\,
            I => \N__20469\
        );

    \I__4853\ : SRMux
    port map (
            O => \N__20670\,
            I => \N__20469\
        );

    \I__4852\ : SRMux
    port map (
            O => \N__20669\,
            I => \N__20469\
        );

    \I__4851\ : SRMux
    port map (
            O => \N__20668\,
            I => \N__20469\
        );

    \I__4850\ : SRMux
    port map (
            O => \N__20667\,
            I => \N__20469\
        );

    \I__4849\ : SRMux
    port map (
            O => \N__20666\,
            I => \N__20469\
        );

    \I__4848\ : SRMux
    port map (
            O => \N__20665\,
            I => \N__20469\
        );

    \I__4847\ : SRMux
    port map (
            O => \N__20664\,
            I => \N__20469\
        );

    \I__4846\ : SRMux
    port map (
            O => \N__20663\,
            I => \N__20469\
        );

    \I__4845\ : SRMux
    port map (
            O => \N__20662\,
            I => \N__20469\
        );

    \I__4844\ : SRMux
    port map (
            O => \N__20661\,
            I => \N__20469\
        );

    \I__4843\ : SRMux
    port map (
            O => \N__20660\,
            I => \N__20469\
        );

    \I__4842\ : SRMux
    port map (
            O => \N__20659\,
            I => \N__20469\
        );

    \I__4841\ : SRMux
    port map (
            O => \N__20658\,
            I => \N__20469\
        );

    \I__4840\ : Glb2LocalMux
    port map (
            O => \N__20655\,
            I => \N__20469\
        );

    \I__4839\ : Glb2LocalMux
    port map (
            O => \N__20652\,
            I => \N__20469\
        );

    \I__4838\ : Glb2LocalMux
    port map (
            O => \N__20649\,
            I => \N__20469\
        );

    \I__4837\ : Glb2LocalMux
    port map (
            O => \N__20646\,
            I => \N__20469\
        );

    \I__4836\ : Glb2LocalMux
    port map (
            O => \N__20643\,
            I => \N__20469\
        );

    \I__4835\ : Glb2LocalMux
    port map (
            O => \N__20640\,
            I => \N__20469\
        );

    \I__4834\ : Glb2LocalMux
    port map (
            O => \N__20637\,
            I => \N__20469\
        );

    \I__4833\ : Glb2LocalMux
    port map (
            O => \N__20634\,
            I => \N__20469\
        );

    \I__4832\ : Glb2LocalMux
    port map (
            O => \N__20631\,
            I => \N__20469\
        );

    \I__4831\ : SRMux
    port map (
            O => \N__20630\,
            I => \N__20469\
        );

    \I__4830\ : SRMux
    port map (
            O => \N__20629\,
            I => \N__20469\
        );

    \I__4829\ : SRMux
    port map (
            O => \N__20628\,
            I => \N__20469\
        );

    \I__4828\ : SRMux
    port map (
            O => \N__20627\,
            I => \N__20469\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__20626\,
            I => \N__20469\
        );

    \I__4826\ : SRMux
    port map (
            O => \N__20625\,
            I => \N__20469\
        );

    \I__4825\ : SRMux
    port map (
            O => \N__20624\,
            I => \N__20469\
        );

    \I__4824\ : SRMux
    port map (
            O => \N__20623\,
            I => \N__20469\
        );

    \I__4823\ : SRMux
    port map (
            O => \N__20622\,
            I => \N__20469\
        );

    \I__4822\ : SRMux
    port map (
            O => \N__20621\,
            I => \N__20469\
        );

    \I__4821\ : SRMux
    port map (
            O => \N__20620\,
            I => \N__20469\
        );

    \I__4820\ : SRMux
    port map (
            O => \N__20619\,
            I => \N__20469\
        );

    \I__4819\ : SRMux
    port map (
            O => \N__20618\,
            I => \N__20469\
        );

    \I__4818\ : SRMux
    port map (
            O => \N__20617\,
            I => \N__20469\
        );

    \I__4817\ : Glb2LocalMux
    port map (
            O => \N__20614\,
            I => \N__20469\
        );

    \I__4816\ : Glb2LocalMux
    port map (
            O => \N__20611\,
            I => \N__20469\
        );

    \I__4815\ : Glb2LocalMux
    port map (
            O => \N__20608\,
            I => \N__20469\
        );

    \I__4814\ : GlobalMux
    port map (
            O => \N__20469\,
            I => \N__20466\
        );

    \I__4813\ : gio2CtrlBuf
    port map (
            O => \N__20466\,
            I => rst_g
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__20463\,
            I => \N__20458\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \N__20454\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20446\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20446\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20439\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20439\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20439\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20433\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20433\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20428\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20428\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \N__20425\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20414\
        );

    \I__4799\ : Span4Mux_s2_v
    port map (
            O => \N__20428\,
            I => \N__20411\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20408\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20391\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20391\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20391\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20391\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20391\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20391\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20391\
        );

    \I__4790\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20391\
        );

    \I__4789\ : Span4Mux_h
    port map (
            O => \N__20414\,
            I => \N__20388\
        );

    \I__4788\ : Sp12to4
    port map (
            O => \N__20411\,
            I => \N__20385\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20408\,
            I => vbuf_tx_data_rdy
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__20391\,
            I => vbuf_tx_data_rdy
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__20388\,
            I => vbuf_tx_data_rdy
        );

    \I__4784\ : Odrv12
    port map (
            O => \N__20385\,
            I => vbuf_tx_data_rdy
        );

    \I__4783\ : CEMux
    port map (
            O => \N__20376\,
            I => \N__20373\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20373\,
            I => \N__20369\
        );

    \I__4781\ : CEMux
    port map (
            O => \N__20372\,
            I => \N__20366\
        );

    \I__4780\ : Span4Mux_s2_v
    port map (
            O => \N__20369\,
            I => \N__20363\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20360\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__20363\,
            I => \N__20357\
        );

    \I__4777\ : Span4Mux_h
    port map (
            O => \N__20360\,
            I => \N__20354\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__20357\,
            I => \N__20351\
        );

    \I__4775\ : Span4Mux_s0_v
    port map (
            O => \N__20354\,
            I => \N__20348\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__20351\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__20348\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__4772\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20337\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \N__20334\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__20341\,
            I => \N__20329\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20326\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20337\,
            I => \N__20323\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20318\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20318\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20313\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20313\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20306\
        );

    \I__4762\ : Span4Mux_s2_h
    port map (
            O => \N__20323\,
            I => \N__20306\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20318\,
            I => \N__20306\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20313\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__20306\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__4758\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20291\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20282\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20282\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20282\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20282\
        );

    \I__4752\ : Span4Mux_s1_v
    port map (
            O => \N__20291\,
            I => \N__20279\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__20282\,
            I => \N__20270\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__20279\,
            I => \N__20267\
        );

    \I__4749\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20256\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20256\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20256\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20256\
        );

    \I__4745\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20256\
        );

    \I__4744\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20253\
        );

    \I__4743\ : Span4Mux_h
    port map (
            O => \N__20270\,
            I => \N__20250\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__20267\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20256\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__20253\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__20250\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__4735\ : Odrv12
    port map (
            O => \N__20232\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20225\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20222\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20219\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20222\,
            I => \Lab_UT.dictrl.N_8_0\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__20219\,
            I => \Lab_UT.dictrl.N_8_0\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20211\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__20208\,
            I => \Lab_UT.dictrl.i8_mux\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20200\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__20204\,
            I => \N__20197\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20193\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20189\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20184\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20184\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20180\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20177\
        );

    \I__4718\ : Span4Mux_s3_v
    port map (
            O => \N__20189\,
            I => \N__20174\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__20184\,
            I => \N__20171\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20168\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__20180\,
            I => bu_rx_data_fast_2
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__20177\,
            I => bu_rx_data_fast_2
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__20174\,
            I => bu_rx_data_fast_2
        );

    \I__4712\ : Odrv12
    port map (
            O => \N__20171\,
            I => bu_rx_data_fast_2
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20168\,
            I => bu_rx_data_fast_2
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__20157\,
            I => \N__20153\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__20156\,
            I => \N__20149\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20144\
        );

    \I__4707\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20144\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20141\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20136\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20132\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__20140\,
            I => \N__20129\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20122\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__20136\,
            I => \N__20119\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20116\
        );

    \I__4699\ : Span4Mux_h
    port map (
            O => \N__20132\,
            I => \N__20113\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20110\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20107\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20104\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20099\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20099\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20096\
        );

    \I__4692\ : Span4Mux_s3_v
    port map (
            O => \N__20119\,
            I => \N__20079\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20079\
        );

    \I__4690\ : Span4Mux_s3_v
    port map (
            O => \N__20113\,
            I => \N__20079\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20079\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20107\,
            I => \N__20079\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20079\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__20099\,
            I => \N__20079\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20096\,
            I => \N__20076\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20071\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20071\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__20079\,
            I => \N__20068\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__20076\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__20071\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__20068\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__20061\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20055\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20055\,
            I => \Lab_UT.dictrl.N_3\
        );

    \I__4675\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20047\
        );

    \I__4674\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20043\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20040\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__20037\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20034\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__20027\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20020\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__20037\,
            I => \N__20020\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20020\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20017\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20014\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20011\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20008\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__20027\,
            I => \N__20003\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__20020\,
            I => \N__20000\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20017\,
            I => \N__19991\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__19991\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__19991\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__19991\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20007\,
            I => \N__19986\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19982\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__19977\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__20000\,
            I => \N__19977\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__19991\,
            I => \N__19974\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19971\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19968\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19965\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19962\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19959\
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__19977\,
            I => bu_rx_data_0
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__19974\,
            I => bu_rx_data_0
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__19971\,
            I => bu_rx_data_0
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19968\,
            I => bu_rx_data_0
        );

    \I__4642\ : Odrv12
    port map (
            O => \N__19965\,
            I => bu_rx_data_0
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19962\,
            I => bu_rx_data_0
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__19959\,
            I => bu_rx_data_0
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__19944\,
            I => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_\
        );

    \I__4638\ : InMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__19938\,
            I => \Lab_UT.dictrl.next_state_RNO_5Z0Z_0\
        );

    \I__4636\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__19932\,
            I => \Lab_UT.dictrl.i9_mux\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__4633\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19911\
        );

    \I__4632\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19911\
        );

    \I__4631\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19906\
        );

    \I__4630\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19903\
        );

    \I__4629\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19900\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19897\
        );

    \I__4627\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19894\
        );

    \I__4626\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19889\
        );

    \I__4625\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19889\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19877\
        );

    \I__4623\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19877\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19874\
        );

    \I__4621\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19869\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19869\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__19906\,
            I => \N__19866\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__19903\,
            I => \N__19860\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19857\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19850\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19850\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__19889\,
            I => \N__19850\
        );

    \I__4613\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19845\
        );

    \I__4612\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19845\
        );

    \I__4611\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19842\
        );

    \I__4610\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19837\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19837\
        );

    \I__4608\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19832\
        );

    \I__4607\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19832\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19822\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__19874\,
            I => \N__19822\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__19869\,
            I => \N__19822\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__19866\,
            I => \N__19822\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19819\
        );

    \I__4601\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19814\
        );

    \I__4600\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19814\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__19860\,
            I => \N__19803\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__19857\,
            I => \N__19803\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__19850\,
            I => \N__19803\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__19845\,
            I => \N__19803\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__19842\,
            I => \N__19803\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__19837\,
            I => \N__19800\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19797\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19831\,
            I => \N__19794\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__19822\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__19819\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__19814\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__19803\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4587\ : Odrv12
    port map (
            O => \N__19800\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__19797\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__19794\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__19779\,
            I => \N__19770\
        );

    \I__4583\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19763\
        );

    \I__4582\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19763\
        );

    \I__4581\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19763\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \N__19760\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__19774\,
            I => \N__19757\
        );

    \I__4578\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19753\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19750\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19763\,
            I => \N__19747\
        );

    \I__4575\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19744\
        );

    \I__4574\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19741\
        );

    \I__4573\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19736\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__19753\,
            I => \N__19733\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19726\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__19747\,
            I => \N__19726\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19726\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19741\,
            I => \N__19723\
        );

    \I__4567\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19720\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19717\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19712\
        );

    \I__4564\ : Span4Mux_s2_v
    port map (
            O => \N__19733\,
            I => \N__19712\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__19726\,
            I => \N__19709\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__19723\,
            I => bu_rx_data_2_rep1
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19720\,
            I => bu_rx_data_2_rep1
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__19717\,
            I => bu_rx_data_2_rep1
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__19712\,
            I => bu_rx_data_2_rep1
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__19709\,
            I => bu_rx_data_2_rep1
        );

    \I__4557\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19692\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19688\
        );

    \I__4555\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19684\
        );

    \I__4554\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19681\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__19692\,
            I => \N__19678\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19675\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__19688\,
            I => \N__19672\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19669\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19663\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19663\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__19678\,
            I => \N__19660\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19653\
        );

    \I__4545\ : Span4Mux_v
    port map (
            O => \N__19672\,
            I => \N__19653\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__19669\,
            I => \N__19653\
        );

    \I__4543\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19650\
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__19663\,
            I => bu_rx_data_0_rep1
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__19660\,
            I => bu_rx_data_0_rep1
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__19653\,
            I => bu_rx_data_0_rep1
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19650\,
            I => bu_rx_data_0_rep1
        );

    \I__4538\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19635\
        );

    \I__4537\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19635\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__19632\,
            I => \Lab_UT.dictrl.N_67_mux\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \N__19623\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \N__19619\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19614\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19611\
        );

    \I__4530\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19608\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__19622\,
            I => \N__19602\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19597\
        );

    \I__4527\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19590\
        );

    \I__4526\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19585\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19585\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19611\,
            I => \N__19582\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__19608\,
            I => \N__19578\
        );

    \I__4522\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19575\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19570\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19570\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19565\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19565\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19562\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19559\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19556\
        );

    \I__4514\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19549\
        );

    \I__4513\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19549\
        );

    \I__4512\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19549\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19542\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19585\,
            I => \N__19542\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__19582\,
            I => \N__19542\
        );

    \I__4508\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19539\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__19578\,
            I => \N__19528\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__19575\,
            I => \N__19528\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__19570\,
            I => \N__19528\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__19565\,
            I => \N__19528\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__19562\,
            I => \N__19528\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__19559\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19556\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__19549\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__19542\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19539\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4497\ : Odrv4
    port map (
            O => \N__19528\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__19515\,
            I => \G_6_0_a6_3_3_cascade_\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19503\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19497\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19491\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19491\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \N__19488\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19485\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19482\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19479\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19472\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19472\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19472\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19468\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19465\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19462\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19455\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__19485\,
            I => \N__19452\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19482\,
            I => \N__19445\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__19479\,
            I => \N__19445\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19445\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19442\
        );

    \I__4475\ : Span4Mux_h
    port map (
            O => \N__19468\,
            I => \N__19435\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19465\,
            I => \N__19435\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__19462\,
            I => \N__19435\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19430\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19430\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19427\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19424\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19455\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__19452\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__19445\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19442\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__19435\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__19430\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19427\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__19424\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19404\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__4458\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19397\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19394\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__19397\,
            I => \N__19388\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__19394\,
            I => \N__19385\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19382\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19377\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19377\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__19388\,
            I => \N__19374\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__19385\,
            I => \N__19371\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__19382\,
            I => bu_rx_data_fast_1
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19377\,
            I => bu_rx_data_fast_1
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__19374\,
            I => bu_rx_data_fast_1
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__19371\,
            I => bu_rx_data_fast_1
        );

    \I__4445\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19352\
        );

    \I__4444\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19352\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19352\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19349\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19342\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19339\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19333\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19333\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19330\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19327\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__19342\,
            I => \N__19322\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__19339\,
            I => \N__19322\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19319\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__19333\,
            I => \N__19316\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__19330\,
            I => bu_rx_data_1_rep1
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19327\,
            I => bu_rx_data_1_rep1
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__19322\,
            I => bu_rx_data_1_rep1
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19319\,
            I => bu_rx_data_1_rep1
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__19316\,
            I => bu_rx_data_1_rep1
        );

    \I__4426\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19301\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19298\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19301\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19298\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__19293\,
            I => \N__19283\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19278\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19275\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19272\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19265\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19265\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19265\
        );

    \I__4415\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19258\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19258\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19258\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__19281\,
            I => \N__19249\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19242\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19242\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19235\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19235\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19258\,
            I => \N__19235\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19232\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__19256\,
            I => \N__19224\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19217\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19217\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19217\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19214\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19211\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19206\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19206\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__19242\,
            I => \N__19201\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__19235\,
            I => \N__19201\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19198\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19231\,
            I => \N__19191\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19191\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19191\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19184\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19184\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19184\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19217\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__19214\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19211\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19206\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__19201\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__19198\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__19191\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19184\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__19167\,
            I => \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__19164\,
            I => \N__19160\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19155\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19155\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19155\,
            I => \Lab_UT.dictrl.N_60\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19143\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19143\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__4371\ : Odrv12
    port map (
            O => \N__19140\,
            I => \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19130\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19127\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19124\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19121\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19117\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19130\,
            I => \N__19114\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19107\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19107\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19107\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19104\
        );

    \I__4360\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19100\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__19114\,
            I => \N__19097\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__19107\,
            I => \N__19094\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19091\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19088\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19100\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__19097\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__19094\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__19091\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__19088\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__19077\,
            I => \G_6_0_a6_2_cascade_\
        );

    \I__4349\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19071\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__19071\,
            I => \Lab_UT.dictrl.G_6_0_0_1\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__19068\,
            I => \Lab_UT.dictrl.G_6_0_0_cascade_\
        );

    \I__4346\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__19059\,
            I => \Lab_UT.dictrl.G_6_0_1_0\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19050\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19050\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__19044\,
            I => \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19037\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19033\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19030\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19024\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__19033\,
            I => \N__19019\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__19030\,
            I => \N__19019\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19029\,
            I => \N__19016\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19011\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19011\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19008\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__19019\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__19016\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19011\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19008\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18993\
        );

    \I__4323\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18993\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__18993\,
            I => \N__18990\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__18990\,
            I => \Lab_UT.dictrl.N_15_0\
        );

    \I__4320\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18983\
        );

    \I__4319\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18978\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18975\
        );

    \I__4317\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18970\
        );

    \I__4316\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18970\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__18978\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__18975\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__18970\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4312\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18957\
        );

    \I__4311\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18957\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__18957\,
            I => \Lab_UT.dictrl.N_59\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__18954\,
            I => \shifter_1_rep1_RNI0FPF_cascade_\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18945\
        );

    \I__4307\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18945\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__18945\,
            I => \Lab_UT.dictrl.N_33_0\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__18942\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__18939\,
            I => \N__18935\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \N__18932\
        );

    \I__4302\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18925\
        );

    \I__4301\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18925\
        );

    \I__4300\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18920\
        );

    \I__4299\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18920\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__18925\,
            I => \Lab_UT.dictrl.G_14_0_1\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__18920\,
            I => \Lab_UT.dictrl.G_14_0_1\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__18915\,
            I => \N__18910\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__18914\,
            I => \N__18907\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__18913\,
            I => \N__18898\
        );

    \I__4293\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18891\
        );

    \I__4292\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18891\
        );

    \I__4291\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18891\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__18905\,
            I => \N__18888\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__18904\,
            I => \N__18883\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__18903\,
            I => \N__18880\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18877\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18872\
        );

    \I__4285\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18872\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__18891\,
            I => \N__18869\
        );

    \I__4283\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18864\
        );

    \I__4282\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18864\
        );

    \I__4281\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18861\
        );

    \I__4280\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18858\
        );

    \I__4279\ : InMux
    port map (
            O => \N__18880\,
            I => \N__18855\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__18877\,
            I => \N__18846\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18846\
        );

    \I__4276\ : Span12Mux_s4_h
    port map (
            O => \N__18869\,
            I => \N__18846\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18864\,
            I => \N__18846\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18861\,
            I => bu_rx_data_3_rep1
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18858\,
            I => bu_rx_data_3_rep1
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__18855\,
            I => bu_rx_data_3_rep1
        );

    \I__4271\ : Odrv12
    port map (
            O => \N__18846\,
            I => bu_rx_data_3_rep1
        );

    \I__4270\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18834\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18834\,
            I => \N__18831\
        );

    \I__4268\ : Odrv12
    port map (
            O => \N__18831\,
            I => \Lab_UT.dictrl.G_14_0_a2_1\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__18828\,
            I => \N_15_cascade_\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__18825\,
            I => \N__18819\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18816\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18807\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18807\
        );

    \I__4262\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18807\
        );

    \I__4261\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18807\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__18807\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__18804\,
            I => \N__18800\
        );

    \I__4258\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18794\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18794\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18791\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18788\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18791\,
            I => \N__18785\
        );

    \I__4253\ : Span4Mux_h
    port map (
            O => \N__18788\,
            I => \N__18782\
        );

    \I__4252\ : Span4Mux_h
    port map (
            O => \N__18785\,
            I => \N__18779\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__18782\,
            I => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__18779\,
            I => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__18774\,
            I => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\
        );

    \I__4248\ : CEMux
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__18765\,
            I => \N__18760\
        );

    \I__4245\ : CEMux
    port map (
            O => \N__18764\,
            I => \N__18757\
        );

    \I__4244\ : CEMux
    port map (
            O => \N__18763\,
            I => \N__18754\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__18760\,
            I => \N__18749\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18749\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18745\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__18749\,
            I => \N__18742\
        );

    \I__4239\ : CEMux
    port map (
            O => \N__18748\,
            I => \N__18739\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__18745\,
            I => \N__18736\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__18742\,
            I => \N__18731\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__18739\,
            I => \N__18731\
        );

    \I__4235\ : Span4Mux_s2_h
    port map (
            O => \N__18736\,
            I => \N__18728\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__18731\,
            I => \N__18725\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__18728\,
            I => \Lab_UT.g0_0\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__18725\,
            I => \Lab_UT.g0_0\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \Lab_UT.dictrl.N_15_0_cascade_\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__18717\,
            I => \Lab_UT.dictrl.N_60_cascade_\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18711\,
            I => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\
        );

    \I__4227\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__18705\,
            I => \N__18701\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18697\
        );

    \I__4224\ : Span4Mux_v
    port map (
            O => \N__18701\,
            I => \N__18694\
        );

    \I__4223\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18691\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18697\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18694\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__18691\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18681\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__4217\ : Span4Mux_h
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__18675\,
            I => \Lab_UT.dictrl.m19_1_0\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18667\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18662\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18662\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18657\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18662\,
            I => \N__18657\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__18657\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18651\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18644\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18644\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__18649\,
            I => \N__18641\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18635\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__18638\,
            I => \N__18630\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__18635\,
            I => \N__18630\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__18630\,
            I => \N__18625\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18622\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18619\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__18625\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18622\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__18619\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__18612\,
            I => \N__18608\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__18611\,
            I => \N__18604\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18593\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18593\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18593\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18593\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18587\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18584\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18579\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18579\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18576\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18573\
        );

    \I__4183\ : Sp12to4
    port map (
            O => \N__18584\,
            I => \N__18568\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__18579\,
            I => \N__18568\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__18576\,
            I => \Lab_UT.next_state_1\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__18573\,
            I => \Lab_UT.next_state_1\
        );

    \I__4179\ : Odrv12
    port map (
            O => \N__18568\,
            I => \Lab_UT.next_state_1\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18554\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18551\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18546\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18551\,
            I => \N__18543\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18538\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18538\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__18546\,
            I => \N__18535\
        );

    \I__4170\ : Span4Mux_v
    port map (
            O => \N__18543\,
            I => \N__18530\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18538\,
            I => \N__18530\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__18535\,
            I => \N__18527\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__18530\,
            I => \N__18524\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__18527\,
            I => \Lab_UT.dictrl.next_state66_2\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18524\,
            I => \Lab_UT.dictrl.next_state66_2\
        );

    \I__4164\ : CEMux
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18511\
        );

    \I__4162\ : CEMux
    port map (
            O => \N__18515\,
            I => \N__18508\
        );

    \I__4161\ : CEMux
    port map (
            O => \N__18514\,
            I => \N__18504\
        );

    \I__4160\ : Span4Mux_s3_h
    port map (
            O => \N__18511\,
            I => \N__18499\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18508\,
            I => \N__18499\
        );

    \I__4158\ : CEMux
    port map (
            O => \N__18507\,
            I => \N__18496\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18504\,
            I => \N__18493\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__18499\,
            I => \N__18488\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18496\,
            I => \N__18488\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__18493\,
            I => \N__18483\
        );

    \I__4153\ : Span4Mux_h
    port map (
            O => \N__18488\,
            I => \N__18483\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__18483\,
            I => \Lab_UT.bu_rx_data_rdy_0\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18474\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__18479\,
            I => \N__18470\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18465\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18477\,
            I => \N__18462\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18474\,
            I => \N__18459\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18456\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18452\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__18469\,
            I => \N__18449\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__18468\,
            I => \N__18446\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18465\,
            I => \N__18442\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__18462\,
            I => \N__18438\
        );

    \I__4140\ : Span4Mux_s3_v
    port map (
            O => \N__18459\,
            I => \N__18433\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18456\,
            I => \N__18433\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18430\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18452\,
            I => \N__18427\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18424\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18413\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18413\
        );

    \I__4133\ : Span4Mux_v
    port map (
            O => \N__18442\,
            I => \N__18410\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18407\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__18438\,
            I => \N__18396\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__18433\,
            I => \N__18396\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18396\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__18427\,
            I => \N__18396\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18396\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18387\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18387\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18387\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18387\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18384\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18381\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18378\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__18410\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__18407\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__18396\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__18387\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18384\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18381\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__18378\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18356\,
            I => \Lab_UT.dictrl.dicRun_1\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18353\,
            I => \Lab_UT.dictrl.dicRun_1\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18342\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18331\
        );

    \I__4105\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18327\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18324\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18321\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18318\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18311\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18311\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18311\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18302\
        );

    \I__4097\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18302\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18302\
        );

    \I__4095\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18302\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18294\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18291\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18288\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__18324\,
            I => \N__18285\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__18321\,
            I => \N__18278\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18278\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18278\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18302\,
            I => \N__18275\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18270\
        );

    \I__4085\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18270\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18263\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18298\,
            I => \N__18263\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18263\
        );

    \I__4081\ : Odrv12
    port map (
            O => \N__18294\,
            I => \Lab_UT.state_2\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18291\,
            I => \Lab_UT.state_2\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__18288\,
            I => \Lab_UT.state_2\
        );

    \I__4078\ : Odrv12
    port map (
            O => \N__18285\,
            I => \Lab_UT.state_2\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__18278\,
            I => \Lab_UT.state_2\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__18275\,
            I => \Lab_UT.state_2\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18270\,
            I => \Lab_UT.state_2\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18263\,
            I => \Lab_UT.state_2\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__18240\,
            I => \N__18236\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18233\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__18236\,
            I => \Lab_UT.LdASones\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18233\,
            I => \Lab_UT.LdASones\
        );

    \I__4067\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18223\
        );

    \I__4066\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18217\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18214\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18211\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18208\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18203\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__18220\,
            I => \N__18198\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18189\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__18214\,
            I => \N__18189\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__18211\,
            I => \N__18184\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18208\,
            I => \N__18184\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18207\,
            I => \N__18181\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18178\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18203\,
            I => \N__18175\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18172\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18167\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18167\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18162\
        );

    \I__4049\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18162\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18159\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18156\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__18189\,
            I => \N__18153\
        );

    \I__4045\ : Span4Mux_h
    port map (
            O => \N__18184\,
            I => \N__18150\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18145\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18178\,
            I => \N__18145\
        );

    \I__4042\ : Span4Mux_v
    port map (
            O => \N__18175\,
            I => \N__18140\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__18172\,
            I => \N__18140\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18167\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18162\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18159\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18156\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__18153\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__18150\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4034\ : Odrv12
    port map (
            O => \N__18145\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__18140\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18107\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18107\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18100\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18100\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18119\,
            I => \N__18100\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18097\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18094\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18087\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18087\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18082\
        );

    \I__4022\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18082\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18074\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__18107\,
            I => \N__18069\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18100\,
            I => \N__18069\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18097\,
            I => \N__18064\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18064\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18061\
        );

    \I__4015\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18058\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18087\,
            I => \N__18053\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18082\,
            I => \N__18053\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18048\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18048\
        );

    \I__4010\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18043\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18043\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18040\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18074\,
            I => \N__18037\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__18069\,
            I => \N__18028\
        );

    \I__4005\ : Span4Mux_v
    port map (
            O => \N__18064\,
            I => \N__18028\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18061\,
            I => \N__18028\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18058\,
            I => \N__18028\
        );

    \I__4002\ : Span4Mux_v
    port map (
            O => \N__18053\,
            I => \N__18025\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__18048\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18043\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18040\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__3998\ : Odrv12
    port map (
            O => \N__18037\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__18028\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__18025\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18012\,
            I => \N__18009\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__18004\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__18008\,
            I => \N__17999\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17994\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__18004\,
            I => \N__17991\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17986\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17986\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17983\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__17998\,
            I => \N__17977\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17972\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17963\
        );

    \I__3984\ : Span4Mux_h
    port map (
            O => \N__17991\,
            I => \N__17963\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__17986\,
            I => \N__17963\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__17983\,
            I => \N__17963\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17958\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17958\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17955\
        );

    \I__3978\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17950\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17950\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17947\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__17972\,
            I => \N__17940\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__17963\,
            I => \N__17940\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__17958\,
            I => \N__17940\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__17955\,
            I => \N__17935\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17950\,
            I => \N__17935\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17947\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__17940\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__17935\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17925\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__17925\,
            I => \N__17922\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__17922\,
            I => \N__17919\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__17919\,
            I => \Lab_UT.dictrl.g1_4_0\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__17916\,
            I => \Lab_UT.dictrl.g1_5_0_cascade_\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__17913\,
            I => \Lab_UT.dictrl.G_14_0_a2_4_2_cascade_\
        );

    \I__3961\ : InMux
    port map (
            O => \N__17910\,
            I => \N__17902\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17902\
        );

    \I__3959\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17897\
        );

    \I__3958\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17897\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__17902\,
            I => \Lab_UT.dictrl.G_14_0_0\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17897\,
            I => \Lab_UT.dictrl.G_14_0_0\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17888\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__17891\,
            I => \N__17885\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17888\,
            I => \N__17878\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17870\
        );

    \I__3951\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17870\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17870\
        );

    \I__3949\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17867\
        );

    \I__3948\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17862\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__17878\,
            I => \N__17859\
        );

    \I__3946\ : InMux
    port map (
            O => \N__17877\,
            I => \N__17856\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17870\,
            I => \N__17853\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17850\
        );

    \I__3943\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17845\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17845\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__17862\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__17859\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__17856\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__17853\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__17850\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17845\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17828\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17824\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17821\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17818\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__17824\,
            I => \N__17815\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__17821\,
            I => \N__17812\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17818\,
            I => \N__17809\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__17815\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__17812\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__17809\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__17802\,
            I => \N__17787\
        );

    \I__3924\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17775\
        );

    \I__3923\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17775\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17775\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17775\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17775\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17766\
        );

    \I__3918\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17766\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17766\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17757\
        );

    \I__3915\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17757\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17791\,
            I => \N__17757\
        );

    \I__3913\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17757\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17752\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17752\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17749\
        );

    \I__3909\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17746\
        );

    \I__3908\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17743\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__17766\,
            I => \N__17740\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17757\,
            I => \N__17733\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__17752\,
            I => \N__17733\
        );

    \I__3904\ : Span4Mux_s3_v
    port map (
            O => \N__17749\,
            I => \N__17733\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17746\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__17743\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__17740\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__17733\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__3898\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17713\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17720\,
            I => \N__17713\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__17719\,
            I => \N__17709\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__17718\,
            I => \N__17705\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__17713\,
            I => \N__17701\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17690\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17690\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17690\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17690\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17690\
        );

    \I__3888\ : Span4Mux_h
    port map (
            O => \N__17701\,
            I => \N__17687\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17690\,
            I => \N__17684\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__17687\,
            I => \Lab_UT.sec2_1\
        );

    \I__3885\ : Odrv12
    port map (
            O => \N__17684\,
            I => \Lab_UT.sec2_1\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17671\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17666\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17666\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__17676\,
            I => \N__17663\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17658\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17658\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17653\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17653\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17650\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17658\,
            I => \N__17647\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__17653\,
            I => \N__17644\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17641\
        );

    \I__3872\ : Span4Mux_v
    port map (
            O => \N__17647\,
            I => \N__17638\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__17644\,
            I => \Lab_UT.LdMtens\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__17641\,
            I => \Lab_UT.LdMtens\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__17638\,
            I => \Lab_UT.LdMtens\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__17631\,
            I => \N__17628\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17625\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17622\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__17622\,
            I => \Lab_UT.didp.countrce4.un13_qPone\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17615\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17612\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__17615\,
            I => \N__17604\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17604\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__17611\,
            I => \N__17600\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17595\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17595\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__17604\,
            I => \N__17592\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17587\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17587\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17595\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__17592\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17587\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17574\,
            I => \Lab_UT.didp.countrce4.q_5_2\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__17571\,
            I => \N__17568\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17565\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17565\,
            I => \N__17562\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__17562\,
            I => \N__17559\
        );

    \I__3844\ : Span4Mux_h
    port map (
            O => \N__17559\,
            I => \N__17555\
        );

    \I__3843\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17552\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__17555\,
            I => \uu0_sec_clkD\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17552\,
            I => \uu0_sec_clkD\
        );

    \I__3840\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17543\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17539\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17543\,
            I => \N__17536\
        );

    \I__3837\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17532\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17529\
        );

    \I__3835\ : Span4Mux_s2_v
    port map (
            O => \N__17536\,
            I => \N__17526\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17523\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__17532\,
            I => \N__17520\
        );

    \I__3832\ : Span4Mux_v
    port map (
            O => \N__17529\,
            I => \N__17513\
        );

    \I__3831\ : Span4Mux_v
    port map (
            O => \N__17526\,
            I => \N__17513\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17523\,
            I => \N__17513\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__17520\,
            I => \N__17507\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__17513\,
            I => \N__17507\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17504\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__17507\,
            I => \N__17501\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17504\,
            I => \o_One_Sec_Pulse\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__17501\,
            I => \o_One_Sec_Pulse\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__17496\,
            I => \N__17488\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__17495\,
            I => \N__17484\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__17494\,
            I => \N__17481\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__17493\,
            I => \N__17477\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17472\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17472\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17465\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17465\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17465\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17462\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__17480\,
            I => \N__17459\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17456\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17449\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17465\,
            I => \N__17449\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17449\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17446\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17443\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__17449\,
            I => \N__17438\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17446\,
            I => \N__17438\
        );

    \I__3804\ : Odrv12
    port map (
            O => \N__17443\,
            I => \oneSecStrb\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__17438\,
            I => \oneSecStrb\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__17433\,
            I => \oneSecStrb_cascade_\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__17430\,
            I => \N__17426\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17423\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17420\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__17423\,
            I => \N__17417\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17414\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__17417\,
            I => \N__17411\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__17414\,
            I => \N__17408\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__17411\,
            I => \Lab_UT.dispString.N_102\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__17408\,
            I => \Lab_UT.dispString.N_102\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17400\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17400\,
            I => \N__17396\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17393\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__17396\,
            I => \N__17390\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17393\,
            I => \N__17387\
        );

    \I__3787\ : Span4Mux_h
    port map (
            O => \N__17390\,
            I => \N__17384\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__17387\,
            I => \N__17381\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__17384\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__17381\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17373\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17373\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__17370\,
            I => \N__17366\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__17369\,
            I => \N__17363\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17366\,
            I => \N__17360\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17355\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__17360\,
            I => \N__17352\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17349\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17346\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17355\,
            I => \N__17343\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__17352\,
            I => \N__17334\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17349\,
            I => \N__17334\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17334\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__17343\,
            I => \N__17334\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__17334\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17325\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17318\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17318\
        );

    \I__3765\ : InMux
    port map (
            O => \N__17328\,
            I => \N__17318\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17325\,
            I => \N__17311\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17318\,
            I => \N__17311\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17306\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17306\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__17311\,
            I => \Lab_UT.LdMones\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17306\,
            I => \Lab_UT.LdMones\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17295\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17289\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17284\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17284\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__17295\,
            I => \N__17281\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17278\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17273\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17273\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17268\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17284\,
            I => \N__17268\
        );

    \I__3748\ : Span4Mux_h
    port map (
            O => \N__17281\,
            I => \N__17265\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17278\,
            I => \N__17262\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__17273\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__17268\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__17265\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3743\ : Odrv12
    port map (
            O => \N__17262\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__17253\,
            I => \N__17249\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__17252\,
            I => \N__17244\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17240\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__17248\,
            I => \N__17235\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__17247\,
            I => \N__17232\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17228\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17243\,
            I => \N__17225\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17222\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17219\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17238\,
            I => \N__17216\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17213\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17208\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17208\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17228\,
            I => \N__17205\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__17225\,
            I => \N__17192\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__17222\,
            I => \N__17192\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17192\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17192\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17192\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__17208\,
            I => \N__17192\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__17205\,
            I => \N__17187\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__17192\,
            I => \N__17187\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__17187\,
            I => \Lab_UT.dictrl.state_i_3_0\
        );

    \I__3719\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17181\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17181\,
            I => \N__17178\
        );

    \I__3717\ : Sp12to4
    port map (
            O => \N__17178\,
            I => \N__17175\
        );

    \I__3716\ : Odrv12
    port map (
            O => \N__17175\,
            I => \Lab_UT.dictrl.state_ret_2_fast\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17169\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17169\,
            I => \N__17165\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__17168\,
            I => \N__17161\
        );

    \I__3712\ : Span4Mux_s3_h
    port map (
            O => \N__17165\,
            I => \N__17158\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17155\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17152\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17158\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17155\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17152\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17142\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__17142\,
            I => \N__17137\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17134\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17131\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__17137\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17134\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17131\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17119\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17114\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17114\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17111\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17114\,
            I => \N__17108\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__17111\,
            I => \Lab_UT.dispString.N_144\
        );

    \I__3693\ : Odrv12
    port map (
            O => \N__17108\,
            I => \Lab_UT.dispString.N_144\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17097\
        );

    \I__3691\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17094\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17091\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17088\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__17097\,
            I => \N__17084\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17078\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17078\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17088\,
            I => \N__17074\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__17087\,
            I => \N__17071\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__17084\,
            I => \N__17068\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17065\
        );

    \I__3681\ : Span4Mux_h
    port map (
            O => \N__17078\,
            I => \N__17062\
        );

    \I__3680\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17059\
        );

    \I__3679\ : Span12Mux_s6_h
    port map (
            O => \N__17074\,
            I => \N__17056\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17053\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__17068\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17065\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__17062\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17059\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3673\ : Odrv12
    port map (
            O => \N__17056\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__17053\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__17040\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17033\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17030\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17033\,
            I => \N__17022\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__17030\,
            I => \N__17019\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17016\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17013\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17008\
        );

    \I__3663\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17008\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17005\
        );

    \I__3661\ : Span4Mux_v
    port map (
            O => \N__17022\,
            I => \N__16998\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__17019\,
            I => \N__16998\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__17016\,
            I => \N__16998\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__17013\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__17008\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__17005\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__16998\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16986\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16986\,
            I => \N__16980\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \N__16975\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16970\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16970\
        );

    \I__3649\ : Span4Mux_v
    port map (
            O => \N__16980\,
            I => \N__16967\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16964\
        );

    \I__3647\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16961\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16958\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__16970\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__16967\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__16964\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16961\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__16958\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3640\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16944\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16944\,
            I => \N__16939\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16936\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16933\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__16939\,
            I => \N__16930\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__16936\,
            I => \N__16927\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16933\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__16930\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__16927\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3631\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__3630\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16914\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__16914\,
            I => \N__16906\
        );

    \I__3628\ : InMux
    port map (
            O => \N__16913\,
            I => \N__16895\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16895\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16895\
        );

    \I__3625\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16895\
        );

    \I__3624\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16895\
        );

    \I__3623\ : Span4Mux_h
    port map (
            O => \N__16906\,
            I => \N__16892\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16895\,
            I => \N__16889\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__16892\,
            I => \Lab_UT.sec2_2\
        );

    \I__3620\ : Odrv12
    port map (
            O => \N__16889\,
            I => \Lab_UT.sec2_2\
        );

    \I__3619\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16875\
        );

    \I__3618\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16868\
        );

    \I__3617\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16868\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16868\
        );

    \I__3615\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16865\
        );

    \I__3614\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16860\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16860\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__16875\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__16868\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__16865\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__16860\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3608\ : InMux
    port map (
            O => \N__16851\,
            I => \N__16848\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16848\,
            I => \N__16845\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__16845\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16839\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16839\,
            I => \N__16835\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16832\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__16835\,
            I => \N__16825\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__16832\,
            I => \N__16825\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16820\
        );

    \I__3599\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16820\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__16825\,
            I => \N__16817\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16814\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__16817\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__3595\ : Odrv12
    port map (
            O => \N__16814\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16805\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16802\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16799\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16802\,
            I => \N__16796\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__16799\,
            I => \N__16793\
        );

    \I__3589\ : Odrv12
    port map (
            O => \N__16796\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__16793\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16785\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__16782\,
            I => \N__16777\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16774\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16771\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__16777\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16774\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16771\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__16764\,
            I => \Lab_UT.didp.countrce3.un13_qPone_cascade_\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__16761\,
            I => \Lab_UT.didp.countrce3.q_5_2_cascade_\
        );

    \I__3577\ : InMux
    port map (
            O => \N__16758\,
            I => \N__16755\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__16755\,
            I => \N__16752\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__16752\,
            I => \Lab_UT.didp.reset_12_1_3\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16749\,
            I => \N__16744\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16738\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16735\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16732\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16743\,
            I => \N__16725\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16725\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16725\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16720\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16735\,
            I => \N__16720\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__16732\,
            I => \N__16717\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16725\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__16720\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__16717\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__16710\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__3560\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16703\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \N__16698\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16703\,
            I => \N__16694\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16691\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16688\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16685\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16682\
        );

    \I__3553\ : Span12Mux_v
    port map (
            O => \N__16694\,
            I => \N__16679\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__16691\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16688\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16685\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__16682\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3548\ : Odrv12
    port map (
            O => \N__16679\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16665\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16665\,
            I => \Lab_UT.didp.countrce3.q_5_3\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16658\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16655\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16658\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16655\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__16650\,
            I => \Lab_UT.didp.un1_dicLdMones_0_cascade_\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16647\,
            I => \N__16644\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__16644\,
            I => \N__16641\
        );

    \I__3538\ : Span4Mux_s1_v
    port map (
            O => \N__16641\,
            I => \N__16638\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__16638\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__3536\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16624\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16624\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16624\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16618\
        );

    \I__3532\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16618\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16613\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16610\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__16618\,
            I => \N__16607\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__16617\,
            I => \N__16604\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16598\
        );

    \I__3526\ : Span4Mux_s1_v
    port map (
            O => \N__16613\,
            I => \N__16595\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16592\
        );

    \I__3524\ : Span4Mux_h
    port map (
            O => \N__16607\,
            I => \N__16589\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16584\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16584\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16581\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16578\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__16598\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__16595\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3517\ : Odrv12
    port map (
            O => \N__16592\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__16589\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16584\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16581\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__16578\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__16560\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16545\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16545\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16545\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16545\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16545\,
            I => \N__16537\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16530\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16530\
        );

    \I__3503\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16530\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16526\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__16540\,
            I => \N__16523\
        );

    \I__3500\ : Span4Mux_s2_v
    port map (
            O => \N__16537\,
            I => \N__16518\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16530\,
            I => \N__16518\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16529\,
            I => \N__16515\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16512\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16509\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__16518\,
            I => \N__16506\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__16515\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__16512\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16509\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__16506\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16494\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16488\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16485\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__16485\,
            I => \uu2.bitmap_pmux_19_ns_1\
        );

    \I__3485\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16476\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16476\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16468\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16457\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16457\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16457\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16457\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16457\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__16468\,
            I => \Lab_UT.sec2_0\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16457\,
            I => \Lab_UT.sec2_0\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__16452\,
            I => \N__16448\
        );

    \I__3474\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16440\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16440\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__16447\,
            I => \N__16437\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__16446\,
            I => \N__16433\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__16445\,
            I => \N__16429\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16426\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16415\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16415\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16415\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16415\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16415\
        );

    \I__3463\ : Span4Mux_s2_v
    port map (
            O => \N__16426\,
            I => \N__16410\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16415\,
            I => \N__16410\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__16410\,
            I => \Lab_UT.sec2_3\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16400\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16393\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16393\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16393\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16390\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16400\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16393\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16390\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16380\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16380\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16374\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__16374\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16367\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16364\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16367\,
            I => \N__16361\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16364\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3444\ : Odrv12
    port map (
            O => \N__16361\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__16356\,
            I => \uu2.N_152_cascade_\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__16353\,
            I => \N__16350\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16344\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16341\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__16348\,
            I => \N__16338\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16335\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__16344\,
            I => \N__16330\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16330\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16327\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16335\,
            I => \N__16324\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__16330\,
            I => \N__16321\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16327\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__16324\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__16321\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16308\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16308\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__16308\,
            I => \N__16305\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__16305\,
            I => \N__16302\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__16302\,
            I => \uu2.bitmap_RNIM5E21Z0Z_314\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16296\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16296\,
            I => \N__16291\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16284\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16284\
        );

    \I__3420\ : Span4Mux_s0_v
    port map (
            O => \N__16291\,
            I => \N__16281\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16276\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16276\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16284\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__16281\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16276\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16269\,
            I => \uu2.un3_w_addr_user_4_cascade_\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16263\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16263\,
            I => \uu2.un3_w_addr_user_5\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16254\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16254\,
            I => \N__16251\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__16251\,
            I => \N__16248\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__16248\,
            I => \uu2.un3_w_addr_user\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16242\,
            I => \N__16239\
        );

    \I__3404\ : Span4Mux_h
    port map (
            O => \N__16239\,
            I => \N__16235\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__16238\,
            I => \N__16228\
        );

    \I__3402\ : Span4Mux_v
    port map (
            O => \N__16235\,
            I => \N__16224\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16217\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16217\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16217\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16210\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16210\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16210\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__16224\,
            I => \N__16207\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16217\,
            I => \N__16204\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16210\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3392\ : Odrv4
    port map (
            O => \N__16207\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__16204\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__16197\,
            I => \uu2.un404_ci_cascade_\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16185\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16182\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16178\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16188\,
            I => \N__16171\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16185\,
            I => \N__16171\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16171\
        );

    \I__3382\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16168\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16178\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__3380\ : Odrv12
    port map (
            O => \N__16171\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16168\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16155\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16155\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16155\,
            I => \N__16150\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16145\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16145\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__16150\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16145\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__16140\,
            I => \N__16136\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16125\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16125\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16125\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16125\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__16125\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16117\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \N__16110\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__16120\,
            I => \N__16107\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__16117\,
            I => \N__16103\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16100\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__16115\,
            I => \N__16095\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16090\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16090\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16085\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16085\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16082\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__16103\,
            I => \N__16077\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16100\,
            I => \N__16077\
        );

    \I__3352\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16072\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16072\
        );

    \I__3350\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16069\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16090\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__16085\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__16082\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__16077\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16072\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__16069\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__16056\,
            I => \N__16053\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16050\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__16050\,
            I => \N__16047\
        );

    \I__3340\ : Span4Mux_h
    port map (
            O => \N__16047\,
            I => \N__16044\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__16044\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16036\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16033\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__16039\,
            I => \N__16030\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16025\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__16033\,
            I => \N__16025\
        );

    \I__3333\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16022\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__16025\,
            I => \uu2.un426_ci_3\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16022\,
            I => \uu2.un426_ci_3\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__16017\,
            I => \N__16013\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16005\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16005\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16005\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16005\,
            I => \N__16002\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__16002\,
            I => \N__15998\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15995\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__15998\,
            I => \uu2.un404_ci\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__15995\,
            I => \uu2.un404_ci\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__15990\,
            I => \N__15987\
        );

    \I__3320\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15984\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15984\,
            I => \N__15981\
        );

    \I__3318\ : Odrv12
    port map (
            O => \N__15981\,
            I => \uu2.vbuf_w_addr_user.un448_ci_0\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15975\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__15975\,
            I => \N__15970\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15965\
        );

    \I__3314\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15965\
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__15970\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__15965\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__3311\ : CEMux
    port map (
            O => \N__15960\,
            I => \N__15957\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__15957\,
            I => \N__15954\
        );

    \I__3309\ : Sp12to4
    port map (
            O => \N__15954\,
            I => \N__15951\
        );

    \I__3308\ : Odrv12
    port map (
            O => \N__15951\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__3307\ : SRMux
    port map (
            O => \N__15948\,
            I => \N__15945\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__15945\,
            I => \N__15942\
        );

    \I__3305\ : Span4Mux_s0_v
    port map (
            O => \N__15942\,
            I => \N__15938\
        );

    \I__3304\ : SRMux
    port map (
            O => \N__15941\,
            I => \N__15935\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__15938\,
            I => \N__15930\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15935\,
            I => \N__15930\
        );

    \I__3301\ : Span4Mux_s0_v
    port map (
            O => \N__15930\,
            I => \N__15926\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15923\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__15926\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_4\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15923\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_4\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15914\
        );

    \I__3296\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15911\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15908\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__15911\,
            I => \N__15905\
        );

    \I__3293\ : Span4Mux_h
    port map (
            O => \N__15908\,
            I => \N__15902\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__15905\,
            I => \N__15899\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__15902\,
            I => \N__15896\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__15899\,
            I => \uu2.N_44\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__15896\,
            I => \uu2.N_44\
        );

    \I__3288\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15882\
        );

    \I__3287\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15882\
        );

    \I__3286\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15882\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__15882\,
            I => \N__15873\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15868\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15868\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15863\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15856\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15856\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15856\
        );

    \I__3278\ : Span4Mux_v
    port map (
            O => \N__15873\,
            I => \N__15853\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15850\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15845\
        );

    \I__3275\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15845\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15863\,
            I => \N__15842\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__15856\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__15853\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__15850\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__15845\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__15842\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15828\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15824\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15821\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15824\,
            I => bu_rx_data_fast_6
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15821\,
            I => bu_rx_data_fast_6
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \N__15812\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15809\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15806\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15809\,
            I => \N__15801\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15806\,
            I => \N__15801\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__15801\,
            I => bu_rx_data_fast_5
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__15798\,
            I => \Lab_UT.dictrl.g1_0_4_cascade_\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15792\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15792\,
            I => \Lab_UT.dictrl.g1_0_xZ0Z1\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15786\,
            I => \Lab_UT.dictrl.g0_5Z0Z_4\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15780\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15780\,
            I => \Lab_UT.dictrl.g0_5_3\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__15777\,
            I => \Lab_UT.dictrl.g1_0_cascade_\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15770\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15767\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15764\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15767\,
            I => \N__15761\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__15764\,
            I => \N__15758\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__15761\,
            I => \N__15755\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__15758\,
            I => \Lab_UT.dictrl.N_55_0\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__15755\,
            I => \Lab_UT.dictrl.N_55_0\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__15750\,
            I => \Lab_UT.dictrl.g0_3_4_cascade_\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15731\
        );

    \I__3239\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15731\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15728\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15744\,
            I => \N__15719\
        );

    \I__3236\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15719\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15719\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15719\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15716\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15711\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15738\,
            I => \N__15711\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15706\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15706\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__15731\,
            I => \N__15699\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15728\,
            I => \N__15699\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15699\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15696\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15691\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__15706\,
            I => \N__15691\
        );

    \I__3222\ : Span4Mux_v
    port map (
            O => \N__15699\,
            I => \N__15688\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__15696\,
            I => bu_rx_data_5
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__15691\,
            I => bu_rx_data_5
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__15688\,
            I => bu_rx_data_5
        );

    \I__3218\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15675\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__15675\,
            I => \N__15672\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__15672\,
            I => \Lab_UT.dictrl.N_72_mux_0\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15662\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15657\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15657\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15652\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15652\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__15662\,
            I => bu_rx_data_6_rep1
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__15657\,
            I => bu_rx_data_6_rep1
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15652\,
            I => bu_rx_data_6_rep1
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \N__15638\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15635\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15630\
        );

    \I__3203\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15630\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15625\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15625\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15635\,
            I => bu_rx_data_7_rep1
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15630\,
            I => bu_rx_data_7_rep1
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__15625\,
            I => bu_rx_data_7_rep1
        );

    \I__3197\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15615\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__15615\,
            I => \Lab_UT.dictrl.g0_3_3\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15604\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15604\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__15610\,
            I => \N__15597\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15593\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15604\,
            I => \N__15590\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15603\,
            I => \N__15584\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15580\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15577\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15574\
        );

    \I__3186\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15571\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15568\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15593\,
            I => \N__15565\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__15590\,
            I => \N__15562\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15559\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15556\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15549\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15549\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15549\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15580\,
            I => bu_rx_data_4
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15577\,
            I => bu_rx_data_4
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__15574\,
            I => bu_rx_data_4
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15571\,
            I => bu_rx_data_4
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15568\,
            I => bu_rx_data_4
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__15565\,
            I => bu_rx_data_4
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__15562\,
            I => bu_rx_data_4
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15559\,
            I => bu_rx_data_4
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15556\,
            I => bu_rx_data_4
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15549\,
            I => bu_rx_data_4
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15516\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15513\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15508\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15508\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__15516\,
            I => \N__15505\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15513\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15508\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__15505\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__15495\,
            I => \N__15491\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15487\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15481\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15481\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15478\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15475\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15481\,
            I => \N__15472\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__15478\,
            I => \N__15469\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15466\
        );

    \I__3147\ : Odrv12
    port map (
            O => \N__15472\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__15469\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15466\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15451\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15451\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15446\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15446\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15451\,
            I => m7_a0
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__15446\,
            I => m7_a0
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__15441\,
            I => \N__15436\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15433\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \N__15430\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15427\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15422\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15422\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15427\,
            I => \N__15419\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__15422\,
            I => \N__15416\
        );

    \I__3130\ : Sp12to4
    port map (
            O => \N__15419\,
            I => \N__15411\
        );

    \I__3129\ : Sp12to4
    port map (
            O => \N__15416\,
            I => \N__15411\
        );

    \I__3128\ : Odrv12
    port map (
            O => \N__15411\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15405\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15405\,
            I => \N__15402\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__15402\,
            I => \N__15395\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15388\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15388\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15388\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15385\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__15395\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__15388\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__15385\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15371\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15371\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__15376\,
            I => \N__15368\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15371\,
            I => \N__15364\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15359\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15359\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__15364\,
            I => bu_rx_data_5_rep1
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__15359\,
            I => bu_rx_data_5_rep1
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__15354\,
            I => \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15348\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15348\,
            I => \N__15345\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__15345\,
            I => \Lab_UT.dictrl.g0_6_3\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__15342\,
            I => \N__15338\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15335\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15332\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__15335\,
            I => \Lab_UT.dictrl.gZ0Z2\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15332\,
            I => \Lab_UT.dictrl.gZ0Z2\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \Lab_UT.dictrl.g0_6_3_cascade_\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15317\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15314\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__15317\,
            I => \Lab_UT.dictrl.g1_1\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15314\,
            I => \Lab_UT.dictrl.g1_1\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15303\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15300\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__15297\,
            I => \Lab_UT.dictrl.N_57_0\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \N_5_cascade_\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15285\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15285\,
            I => \Lab_UT.dictrl.N_59_1_0\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15276\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15276\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15276\,
            I => \Lab_UT.dictrl.i8_mux_0\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15270\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15270\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__15267\,
            I => \Lab_UT.dictrl.m22_xZ0Z1_cascade_\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15259\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15253\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15253\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15259\,
            I => \N__15250\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15247\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__15253\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__15250\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15247\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__15240\,
            I => \Lab_UT.dictrl.N_72_mux_cascade_\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15234\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__15234\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \Lab_UT.dictrl.m34_0_cascade_\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__15228\,
            I => \Lab_UT.dictrl.next_state_1_3_cascade_\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__15225\,
            I => \N__15221\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15217\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15210\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15210\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15217\,
            I => \N__15210\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15210\,
            I => \N__15207\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__15207\,
            I => \N__15204\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__15204\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15201\,
            I => \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15186\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15186\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15186\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15186\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15186\,
            I => \N__15183\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__15183\,
            I => \Lab_UT.dictrl.N_26_0\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15177\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15177\,
            I => \Lab_UT.dictrl.m34_0\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15174\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15168\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15168\,
            I => \Lab_UT.dictrl.N_60_0_0\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15159\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15159\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15159\,
            I => \N__15156\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__15156\,
            I => \Lab_UT.dictrl.m19_1\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15149\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15146\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15149\,
            I => \N__15141\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15146\,
            I => \N__15141\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__15141\,
            I => \Lab_UT.dictrl.N_22\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__15138\,
            I => \N__15135\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15132\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15132\,
            I => \N__15129\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__15129\,
            I => \Lab_UT.dictrl.next_state_0_1\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \N__15123\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15120\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__15120\,
            I => \N__15117\
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__15117\,
            I => \Lab_UT.dictrl.g2_0_0\
        );

    \I__3029\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15104\
        );

    \I__3028\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15104\
        );

    \I__3027\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15104\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__15111\,
            I => \N__15101\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__15104\,
            I => \N__15098\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15095\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__15098\,
            I => \Lab_UT.dictrl.state_i_4_2\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15095\,
            I => \Lab_UT.dictrl.state_i_4_2\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__15090\,
            I => \Lab_UT.dictrl.N_20_0_0_cascade_\
        );

    \I__3020\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15084\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__15084\,
            I => \N__15081\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__15081\,
            I => \N__15078\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__15078\,
            I => \Lab_UT.dictrl.N_22_0_0\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15064\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15064\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15060\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15051\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15051\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15051\
        );

    \I__3010\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15051\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15064\,
            I => \N__15048\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15045\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15060\,
            I => \Lab_UT.next_state_0\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__15051\,
            I => \Lab_UT.next_state_0\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__15048\,
            I => \Lab_UT.next_state_0\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15045\,
            I => \Lab_UT.next_state_0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15036\,
            I => \Lab_UT.next_state_1_0_0_1_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15024\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15015\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15015\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15015\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15029\,
            I => \N__15015\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15010\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15010\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__15024\,
            I => \N__15007\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15015\,
            I => \Lab_UT.next_state_2\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15010\,
            I => \Lab_UT.next_state_2\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__15007\,
            I => \Lab_UT.next_state_2\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14987\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14987\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14987\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14987\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14984\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__14987\,
            I => \N__14981\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14975\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__14981\,
            I => \N__14971\
        );

    \I__2983\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14968\
        );

    \I__2982\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14963\
        );

    \I__2981\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14963\
        );

    \I__2980\ : Sp12to4
    port map (
            O => \N__14975\,
            I => \N__14958\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14955\
        );

    \I__2978\ : Sp12to4
    port map (
            O => \N__14971\,
            I => \N__14948\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__14968\,
            I => \N__14948\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14963\,
            I => \N__14948\
        );

    \I__2975\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14945\
        );

    \I__2974\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14942\
        );

    \I__2973\ : Span12Mux_s4_v
    port map (
            O => \N__14958\,
            I => \N__14937\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14937\
        );

    \I__2971\ : Span12Mux_s11_h
    port map (
            O => \N__14948\,
            I => \N__14934\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__14945\,
            I => bu_rx_data_rdy
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__14942\,
            I => bu_rx_data_rdy
        );

    \I__2968\ : Odrv12
    port map (
            O => \N__14937\,
            I => bu_rx_data_rdy
        );

    \I__2967\ : Odrv12
    port map (
            O => \N__14934\,
            I => bu_rx_data_rdy
        );

    \I__2966\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14922\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__14922\,
            I => \Lab_UT.didp.g0_0_2Z0Z_1\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__14919\,
            I => \N__14916\
        );

    \I__2963\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14911\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__14915\,
            I => \N__14907\
        );

    \I__2961\ : IoInMux
    port map (
            O => \N__14914\,
            I => \N__14904\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14911\,
            I => \N__14901\
        );

    \I__2959\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14898\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14895\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__14904\,
            I => \N__14892\
        );

    \I__2956\ : Sp12to4
    port map (
            O => \N__14901\,
            I => \N__14885\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__14898\,
            I => \N__14885\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14885\
        );

    \I__2953\ : Span4Mux_s0_h
    port map (
            O => \N__14892\,
            I => \N__14882\
        );

    \I__2952\ : Odrv12
    port map (
            O => \N__14885\,
            I => rst
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__14882\,
            I => rst
        );

    \I__2950\ : InMux
    port map (
            O => \N__14877\,
            I => \N__14874\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__14874\,
            I => \Lab_UT.didp.g0_0Z0Z_2\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14865\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14865\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__14865\,
            I => \N__14862\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__14862\,
            I => \N__14859\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__14859\,
            I => \Lab_UT.dictrl.next_state6\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__14856\,
            I => \Lab_UT.dictrl.N_20_cascade_\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__14853\,
            I => \Lab_UT.dictrl.un15_loadalarm_0_cascade_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14847\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__14847\,
            I => \Lab_UT.dictrl.loadalarm_0_0\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14840\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14837\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14840\,
            I => \N__14834\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__14837\,
            I => \N__14831\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__14834\,
            I => \Lab_UT.LdAStens\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__14831\,
            I => \Lab_UT.LdAStens\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__14826\,
            I => \N__14823\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14819\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14816\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14819\,
            I => \Lab_UT.dictrl.dicLdAMones_1\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14816\,
            I => \Lab_UT.dictrl.dicLdAMones_1\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__14808\,
            I => \N__14805\
        );

    \I__2926\ : Span4Mux_h
    port map (
            O => \N__14805\,
            I => \N__14802\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__14802\,
            I => \Lab_UT.LdAMones\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__14799\,
            I => \Lab_UT.LdAMones_cascade_\
        );

    \I__2923\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14793\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14793\,
            I => \Lab_UT.dictrl.g0_1_mb_rn_0\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__14790\,
            I => \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14784\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__14784\,
            I => \N__14780\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14777\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__14780\,
            I => \N__14774\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__14777\,
            I => \N__14771\
        );

    \I__2915\ : Span4Mux_v
    port map (
            O => \N__14774\,
            I => \N__14768\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__14771\,
            I => \N__14765\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__14768\,
            I => \Lab_UT.dictrl.N_57_1\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__14765\,
            I => \Lab_UT.dictrl.N_57_1\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__14760\,
            I => \N__14757\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14754\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14754\,
            I => \N__14750\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__14753\,
            I => \N__14747\
        );

    \I__2907\ : Span4Mux_s2_v
    port map (
            O => \N__14750\,
            I => \N__14744\
        );

    \I__2906\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14741\
        );

    \I__2905\ : Span4Mux_v
    port map (
            O => \N__14744\,
            I => \N__14738\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14735\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__14738\,
            I => \N__14732\
        );

    \I__2902\ : Span4Mux_h
    port map (
            O => \N__14735\,
            I => \N__14729\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__14732\,
            I => \Lab_UT.dictrl.N_55_1\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__14729\,
            I => \Lab_UT.dictrl.N_55_1\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14721\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14721\,
            I => \N__14717\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__14720\,
            I => \N__14713\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__14717\,
            I => \N__14710\
        );

    \I__2895\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14705\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14705\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__14710\,
            I => \N__14702\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14699\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__14702\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__2890\ : Odrv12
    port map (
            O => \N__14699\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__14694\,
            I => \Lab_UT.dictrl.next_state_1_2_cascade_\
        );

    \I__2888\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14685\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14685\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14685\,
            I => \Lab_UT.dictrl.g0_1_mb_sn\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14675\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14675\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14672\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14675\,
            I => \N__14669\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__14672\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2880\ : Odrv12
    port map (
            O => \N__14669\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14661\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14661\,
            I => \N__14652\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14639\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14639\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14639\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14639\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14639\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14639\
        );

    \I__2871\ : Span4Mux_s2_v
    port map (
            O => \N__14652\,
            I => \N__14636\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14639\,
            I => \N__14633\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__14636\,
            I => \Lab_UT.min1_2\
        );

    \I__2868\ : Odrv12
    port map (
            O => \N__14633\,
            I => \Lab_UT.min1_2\
        );

    \I__2867\ : CEMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14625\,
            I => \N__14622\
        );

    \I__2865\ : Span4Mux_v
    port map (
            O => \N__14622\,
            I => \N__14618\
        );

    \I__2864\ : CEMux
    port map (
            O => \N__14621\,
            I => \N__14615\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__14618\,
            I => \N__14612\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14615\,
            I => \N__14609\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__14612\,
            I => \Lab_UT.didp.regrce3.LdAMones_0\
        );

    \I__2860\ : Odrv12
    port map (
            O => \N__14609\,
            I => \Lab_UT.didp.regrce3.LdAMones_0\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14595\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14595\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14595\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__14595\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14588\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14585\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__14588\,
            I => \N__14580\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14585\,
            I => \N__14580\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__14580\,
            I => \N__14576\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14573\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__14576\,
            I => \N__14570\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14567\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__14570\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2846\ : Odrv12
    port map (
            O => \N__14567\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__14562\,
            I => \Lab_UT.dispString.N_118_cascade_\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14559\,
            I => \N__14556\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__14550\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_1\
        );

    \I__2840\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14543\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__14546\,
            I => \N__14540\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__14543\,
            I => \N__14537\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14534\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__14537\,
            I => \N__14528\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14534\,
            I => \N__14528\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14525\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__14528\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14525\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14516\
        );

    \I__2830\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14512\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14509\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14506\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14501\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__14509\,
            I => \N__14501\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14506\,
            I => \N__14498\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__14501\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__14498\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__14493\,
            I => \N__14487\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__14492\,
            I => \N__14483\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__14491\,
            I => \N__14479\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14490\,
            I => \N__14475\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14462\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14462\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14462\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14462\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14462\
        );

    \I__2813\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14462\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__14475\,
            I => \N__14457\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14457\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__14457\,
            I => \Lab_UT.min1_1\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14443\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14443\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14443\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14440\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14450\,
            I => \N__14436\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__14443\,
            I => \N__14431\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14431\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14439\,
            I => \N__14426\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14426\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__14431\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14426\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14417\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14414\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__14417\,
            I => \N__14411\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14414\,
            I => \N__14405\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__14411\,
            I => \N__14405\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14402\
        );

    \I__2792\ : Span4Mux_v
    port map (
            O => \N__14405\,
            I => \N__14399\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14402\,
            I => \N__14396\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__14399\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__14396\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14391\,
            I => \N__14373\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14373\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14373\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14388\,
            I => \N__14373\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14373\
        );

    \I__2783\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14373\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__14373\,
            I => \N__14369\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14366\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__14369\,
            I => \Lab_UT.sec1_2\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14366\,
            I => \Lab_UT.sec1_2\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14357\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14352\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14348\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14343\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14355\,
            I => \N__14340\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__14352\,
            I => \N__14337\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14333\
        );

    \I__2771\ : Span4Mux_h
    port map (
            O => \N__14348\,
            I => \N__14330\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14327\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14324\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__14343\,
            I => \N__14317\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14317\
        );

    \I__2766\ : Span4Mux_s2_v
    port map (
            O => \N__14337\,
            I => \N__14317\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14314\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__14333\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__14330\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14327\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__14324\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__14317\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__14314\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14298\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14295\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__14295\,
            I => \N__14289\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__14294\,
            I => \N__14286\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14283\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14280\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__14289\,
            I => \N__14277\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14286\,
            I => \N__14274\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14283\,
            I => \N__14271\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14280\,
            I => \Lab_UT.LdSones\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__14277\,
            I => \Lab_UT.LdSones\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14274\,
            I => \Lab_UT.LdSones\
        );

    \I__2746\ : Odrv12
    port map (
            O => \N__14271\,
            I => \Lab_UT.LdSones\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14262\,
            I => \Lab_UT.didp.countrce1.un13_qPone_cascade_\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__14259\,
            I => \N__14255\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14258\,
            I => \N__14252\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14246\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14246\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14243\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14246\,
            I => \N__14239\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14243\,
            I => \N__14236\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14233\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__14239\,
            I => \N__14230\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__14236\,
            I => \N__14227\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14224\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__14230\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__14227\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__2731\ : Odrv12
    port map (
            O => \N__14224\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__14217\,
            I => \Lab_UT.didp.countrce1.q_5_2_cascade_\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14211\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14211\,
            I => \N__14205\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14202\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14199\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14196\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__14205\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14202\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14199\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14196\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14178\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14178\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14178\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14175\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__14175\,
            I => \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14169\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14169\,
            I => \N__14166\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__14166\,
            I => \N__14163\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__14163\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14160\,
            I => \N__14155\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__14159\,
            I => \N__14152\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14140\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14155\,
            I => \N__14140\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14140\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14140\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__14150\,
            I => \N__14137\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \N__14134\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14130\
        );

    \I__2702\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14123\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14123\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14133\,
            I => \N__14123\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__14130\,
            I => \N__14118\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__14123\,
            I => \N__14118\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__14118\,
            I => \Lab_UT.min2_1\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14115\,
            I => \N__14106\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__14114\,
            I => \N__14103\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14100\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__14112\,
            I => \N__14097\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14094\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__14110\,
            I => \N__14091\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__14109\,
            I => \N__14088\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14085\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14076\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14076\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14076\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14076\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14071\
        );

    \I__2683\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14071\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__14085\,
            I => \Lab_UT.sec1_3\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__14076\,
            I => \Lab_UT.sec1_3\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14071\,
            I => \Lab_UT.sec1_3\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14055\
        );

    \I__2678\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14042\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14042\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14042\
        );

    \I__2675\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14042\
        );

    \I__2674\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14042\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14042\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__14055\,
            I => \Lab_UT.sec1_0\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14042\,
            I => \Lab_UT.sec1_0\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14034\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__14034\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14028\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__14028\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14022\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14022\,
            I => \uu2.bitmap_pmux_17_ns_1\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__14019\,
            I => \N__14014\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__14018\,
            I => \N__14011\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14004\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14004\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14004\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14004\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13998\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__13998\,
            I => \N__13995\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__13995\,
            I => \N__13992\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__13992\,
            I => \uu2.bitmap_pmux_16_ns_1\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13989\,
            I => \N__13986\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13986\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13980\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13980\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__2650\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13965\
        );

    \I__2649\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13965\
        );

    \I__2648\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13965\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13965\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__13965\,
            I => \N__13959\
        );

    \I__2645\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13952\
        );

    \I__2644\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13952\
        );

    \I__2643\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13952\
        );

    \I__2642\ : Odrv12
    port map (
            O => \N__13959\,
            I => \Lab_UT.min2_0\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__13952\,
            I => \Lab_UT.min2_0\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__13947\,
            I => \N__13942\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__13946\,
            I => \N__13937\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__13945\,
            I => \N__13932\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13942\,
            I => \N__13923\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13941\,
            I => \N__13923\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13923\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13923\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13916\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13916\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13916\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13923\,
            I => \Lab_UT.min2_3\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__13916\,
            I => \Lab_UT.min2_3\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13899\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13899\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13899\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13899\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__13899\,
            I => \N__13893\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13886\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13886\
        );

    \I__2621\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13886\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__13893\,
            I => \Lab_UT.min2_2\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13886\,
            I => \Lab_UT.min2_2\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13878\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__13878\,
            I => \N__13875\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__13875\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13866\
        );

    \I__2614\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13858\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13858\
        );

    \I__2612\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13858\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__13866\,
            I => \N__13855\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13850\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13858\,
            I => \N__13845\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__13855\,
            I => \N__13845\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13840\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13840\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__13850\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__13845\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13840\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2602\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13818\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13818\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13818\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13818\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13813\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13813\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13810\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__13818\,
            I => \Lab_UT.sec1_1\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__13813\,
            I => \Lab_UT.sec1_1\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13810\,
            I => \Lab_UT.sec1_1\
        );

    \I__2592\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13800\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__13800\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13794\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__13794\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__13791\,
            I => \N__13786\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \N__13783\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__13789\,
            I => \N__13779\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13774\
        );

    \I__2584\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13771\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13766\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13766\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13761\
        );

    \I__2580\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13761\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13774\,
            I => \N__13758\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13771\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__13766\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13761\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__13758\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2574\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13746\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__13746\,
            I => \uu2.bitmap_pmux_26_bm_1\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13740\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13740\,
            I => \N__13737\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__13737\,
            I => \uu2.bitmap_RNIP2JO1Z0Z_34\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13734\,
            I => \N__13731\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__13731\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13722\
        );

    \I__2566\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13714\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13714\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13714\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__13722\,
            I => \N__13711\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__13721\,
            I => \N__13706\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13714\,
            I => \N__13703\
        );

    \I__2560\ : Span12Mux_s6_v
    port map (
            O => \N__13711\,
            I => \N__13700\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13693\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13693\
        );

    \I__2557\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13693\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__13703\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__13700\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13693\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__13686\,
            I => \N__13683\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13679\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13676\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__13679\,
            I => \N__13672\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13676\,
            I => \N__13669\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13666\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__13672\,
            I => \N__13663\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__13669\,
            I => \N__13660\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__13666\,
            I => \N__13657\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__13663\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__13660\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__13657\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13650\,
            I => \N__13646\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13649\,
            I => \N__13643\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13640\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13643\,
            I => \N__13637\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__13640\,
            I => \N__13632\
        );

    \I__2536\ : Span4Mux_s2_v
    port map (
            O => \N__13637\,
            I => \N__13632\
        );

    \I__2535\ : Span4Mux_v
    port map (
            O => \N__13632\,
            I => \N__13628\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13625\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__13628\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13625\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13616\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13613\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13609\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13613\,
            I => \N__13606\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13603\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__13609\,
            I => \N__13600\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__13606\,
            I => \N__13597\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13603\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__13600\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__13597\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13586\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13583\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13580\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13576\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__13580\,
            I => \N__13573\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13570\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__13576\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__13573\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13570\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13554\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13541\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13541\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13541\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13541\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13541\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13541\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13554\,
            I => \Lab_UT.min1_0\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13541\,
            I => \Lab_UT.min1_0\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13531\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13526\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13526\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13531\,
            I => \N__13523\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13520\
        );

    \I__2498\ : Span4Mux_h
    port map (
            O => \N__13523\,
            I => \N__13517\
        );

    \I__2497\ : Span4Mux_h
    port map (
            O => \N__13520\,
            I => \N__13514\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__13517\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__13514\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13505\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13502\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13505\,
            I => \N__13499\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13502\,
            I => \N__13492\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__13499\,
            I => \N__13492\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13486\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13486\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__13492\,
            I => \N__13483\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13480\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13486\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__13483\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13480\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__13473\,
            I => \N__13470\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13464\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \N__13460\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__13468\,
            I => \N__13456\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__13467\,
            I => \N__13452\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13464\,
            I => \N__13449\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13436\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13436\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13436\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13436\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13455\,
            I => \N__13436\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13436\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__13449\,
            I => \Lab_UT.min1_3\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__13436\,
            I => \Lab_UT.min1_3\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__13431\,
            I => \N__13428\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13428\,
            I => \N__13423\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__13427\,
            I => \N__13419\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__13426\,
            I => \N__13414\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13423\,
            I => \N__13410\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13397\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13419\,
            I => \N__13397\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13397\
        );

    \I__2460\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13397\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13397\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13397\
        );

    \I__2457\ : Span4Mux_s2_v
    port map (
            O => \N__13410\,
            I => \N__13394\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N__13391\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__13394\,
            I => \uu2.N_37\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__13391\,
            I => \uu2.N_37\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13377\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13377\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13374\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13366\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13363\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13377\,
            I => \N__13360\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13374\,
            I => \N__13357\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13350\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13372\,
            I => \N__13350\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13350\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13345\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13345\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13366\,
            I => \N__13342\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13363\,
            I => \N__13339\
        );

    \I__2439\ : Span4Mux_h
    port map (
            O => \N__13360\,
            I => \N__13336\
        );

    \I__2438\ : Odrv12
    port map (
            O => \N__13357\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13350\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__13345\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__13342\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__13339\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__13336\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__13323\,
            I => \N__13320\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13317\,
            I => \uu2.N_45\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__13308\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__13305\,
            I => \N__13301\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13298\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13290\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13287\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13282\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13282\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13295\,
            I => \N__13275\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13275\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13275\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13290\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2416\ : Odrv12
    port map (
            O => \N__13287\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__13282\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__13275\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13257\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13257\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13253\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13250\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13246\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13243\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__13256\,
            I => \N__13237\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13234\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13231\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13228\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13246\,
            I => \N__13225\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__13243\,
            I => \N__13222\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13242\,
            I => \N__13213\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13213\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13240\,
            I => \N__13213\
        );

    \I__2398\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13213\
        );

    \I__2397\ : Span4Mux_h
    port map (
            O => \N__13234\,
            I => \N__13208\
        );

    \I__2396\ : Span4Mux_h
    port map (
            O => \N__13231\,
            I => \N__13208\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13228\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__13225\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__13222\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13213\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__13208\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13197\,
            I => \N__13194\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13194\,
            I => \N__13190\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__13193\,
            I => \N__13185\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__13190\,
            I => \N__13180\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13189\,
            I => \N__13173\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13173\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13173\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13168\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13168\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__13180\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13173\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13168\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13158\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13158\,
            I => \N__13155\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__13155\,
            I => \N__13152\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__13152\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13149\,
            I => \N__13146\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13146\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13140\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13140\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13134\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__13134\,
            I => \uu2.bitmap_pmux_20_ns_1\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13128\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__13125\,
            I => \Lab_UT.dictrl.g1_1_4_cascade_\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13119\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__13116\,
            I => \Lab_UT.dictrl.g1_1Z0Z_5\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__13113\,
            I => \N__13108\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \N__13105\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13094\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13094\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13084\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13084\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13084\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13081\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13078\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13073\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13073\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13070\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13065\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13065\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13062\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13059\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13054\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13054\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13049\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__13070\,
            I => \N__13049\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__13065\,
            I => \N__13042\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13062\,
            I => \N__13042\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__13059\,
            I => \N__13042\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__13054\,
            I => bu_rx_data_7
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__13049\,
            I => bu_rx_data_7
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__13042\,
            I => bu_rx_data_7
        );

    \I__2336\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13029\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13034\,
            I => \N__13029\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13029\,
            I => \N__13025\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13028\,
            I => \N__13022\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__13025\,
            I => \N__13017\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13022\,
            I => \N__13017\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__13017\,
            I => \N__13013\
        );

    \I__2329\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13010\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__13013\,
            I => \N__13005\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__13010\,
            I => \N__13005\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__13005\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12996\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12996\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12996\,
            I => bu_rx_data_fast_7
        );

    \I__2322\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12983\
        );

    \I__2321\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12983\
        );

    \I__2320\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12983\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__12990\,
            I => \N__12978\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__12983\,
            I => \N__12975\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12982\,
            I => \N__12968\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12968\
        );

    \I__2315\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12968\
        );

    \I__2314\ : Span4Mux_h
    port map (
            O => \N__12975\,
            I => \N__12965\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__12968\,
            I => \uu2.N_40\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__12965\,
            I => \uu2.N_40\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__12960\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__12957\,
            I => \Lab_UT.dictrl.m22Z0Z_1_cascade_\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12951\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12951\,
            I => \Lab_UT.dictrl.N_72_mux_1\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__12948\,
            I => \N__12945\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12942\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__12942\,
            I => \Lab_UT.dictrl.g1_1_0_0\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12935\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12932\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__12935\,
            I => \N__12929\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__12932\,
            I => \Lab_UT.dictrl.m22Z0Z_1\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__12929\,
            I => \Lab_UT.dictrl.m22Z0Z_1\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12921\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__12921\,
            I => \Lab_UT.dictrl.g1_1_0\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \N__12915\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12912\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__12912\,
            I => \N__12909\
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__12909\,
            I => \Lab_UT.dictrl.g1_rn_0\
        );

    \I__2293\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12903\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12903\,
            I => \N__12900\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__12900\,
            I => \N__12896\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12893\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__12896\,
            I => \Lab_UT.dictrl.m34Z0Z_1\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12893\,
            I => \Lab_UT.dictrl.m34Z0Z_1\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__12888\,
            I => \N__12884\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__12887\,
            I => \N__12881\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12878\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12875\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__12878\,
            I => bu_rx_data_fast_3
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__12875\,
            I => bu_rx_data_fast_3
        );

    \I__2281\ : InMux
    port map (
            O => \N__12870\,
            I => \N__12864\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12864\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12864\,
            I => \N__12861\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__12861\,
            I => bu_rx_data_fast_0
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__12858\,
            I => \Lab_UT.dictrl.m13_out_cascade_\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__12855\,
            I => \Lab_UT.dictrl.N_18_0_0_cascade_\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12849\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12849\,
            I => \Lab_UT.dictrl.G_25_i_o3_5\
        );

    \I__2273\ : InMux
    port map (
            O => \N__12846\,
            I => \N__12843\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12843\,
            I => \N__12840\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__12840\,
            I => \Lab_UT.dictrl.G_25_i_o3_4\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__12837\,
            I => \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12831\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12831\,
            I => \Lab_UT.dictrl.N_11\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__12828\,
            I => \Lab_UT.dictrl.m34Z0Z_1_cascade_\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12818\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12813\
        );

    \I__2264\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12813\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12801\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12801\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12818\,
            I => \N__12798\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12795\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12790\
        );

    \I__2258\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12790\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12785\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12785\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12778\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12778\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12778\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12801\,
            I => bu_rx_data_6
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__12798\,
            I => bu_rx_data_6
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__12795\,
            I => bu_rx_data_6
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__12790\,
            I => bu_rx_data_6
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__12785\,
            I => bu_rx_data_6
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12778\,
            I => bu_rx_data_6
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__12765\,
            I => \Lab_UT.i8_mux_0_cascade_\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \N__12759\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12756\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12756\,
            I => \Lab_UT.dictrl.g0_0_sn\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__12753\,
            I => \Lab_UT.dictrl.g1_1_0_1_cascade_\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12747\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__12747\,
            I => \Lab_UT.g1\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__12741\,
            I => \Lab_UT.dictrl.g0_0_rn_0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__12732\,
            I => \Lab_UT.dictrl.G_25_i_0\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__12726\,
            I => \Lab_UT.dictrl.G_25_i_1\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12720\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12717\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__12717\,
            I => \Lab_UT.dictrl.g2Z0Z_0\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__12714\,
            I => \N__12711\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12708\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12708\,
            I => \Lab_UT.dictrl.g0_6_3_0\
        );

    \I__2226\ : CEMux
    port map (
            O => \N__12705\,
            I => \N__12702\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12702\,
            I => \N__12699\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__12699\,
            I => \N__12696\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__12696\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__12693\,
            I => \Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__12690\,
            I => \Lab_UT.dictrl.G_25_i_a5_1_0_cascade_\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12684\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12684\,
            I => \N__12681\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__12681\,
            I => \N__12678\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__12678\,
            I => \Lab_UT.didp.N_90\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12672\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__12672\,
            I => \Lab_UT.LdSones_i_4\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12666\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12666\,
            I => \N__12663\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__12660\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12648\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12648\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12648\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__12648\,
            I => \N__12642\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12637\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12637\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12634\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__12642\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__12637\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12634\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__12627\,
            I => \N__12621\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__12626\,
            I => \N__12617\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__12625\,
            I => \N__12612\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__12624\,
            I => \N__12609\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12604\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12604\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12601\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12598\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12591\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12591\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12591\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12586\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12586\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12598\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__12591\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__12586\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__12579\,
            I => \N__12576\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12573\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__12573\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12567\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__12567\,
            I => \Lab_UT.didp.countrce1.q_5_1\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12560\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__12563\,
            I => \N__12555\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12560\,
            I => \N__12552\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12549\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12546\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12543\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__12552\,
            I => \N__12539\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12549\,
            I => \N__12532\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12532\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12543\,
            I => \N__12532\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12529\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__12539\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__12532\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12529\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12519\,
            I => \N__12514\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12518\,
            I => \N__12511\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12508\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__12514\,
            I => \N__12503\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12511\,
            I => \N__12503\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12508\,
            I => \N__12500\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__12503\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__12500\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12492\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__2154\ : Span4Mux_h
    port map (
            O => \N__12489\,
            I => \N__12486\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__12486\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_0\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12477\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12477\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12477\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12471\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__12468\,
            I => \Lab_UT.didp.un1_dicLdStens_0_cascade_\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__12465\,
            I => \N__12460\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12454\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12454\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12449\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12449\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12454\,
            I => \N__12446\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12443\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__12446\,
            I => \N__12440\
        );

    \I__2138\ : Span4Mux_h
    port map (
            O => \N__12443\,
            I => \N__12437\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__12440\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__12437\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12426\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12426\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12426\,
            I => \N__12423\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__12423\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12417\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12417\,
            I => \N__12414\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__12414\,
            I => \N__12411\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__12411\,
            I => \Lab_UT.didp.countrce1.q_5_0\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12405\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12405\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12398\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12394\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__12398\,
            I => \N__12391\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12388\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12394\,
            I => \N__12385\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__12391\,
            I => \N__12382\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12388\,
            I => \N__12379\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__12385\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__12382\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2116\ : Odrv12
    port map (
            O => \N__12379\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__12366\,
            I => \N__12361\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12356\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12356\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__12361\,
            I => \N__12353\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12356\,
            I => \N__12350\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__12353\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__12350\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__12345\,
            I => \N__12342\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12339\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__12339\,
            I => \Lab_UT.didp.countrce2.N_93\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12333\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12333\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__12330\,
            I => \Lab_UT.didp.countrce2.N_96_cascade_\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12324\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__12324\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12315\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__12312\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__12309\,
            I => \N__12302\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12299\
        );

    \I__2092\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12296\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12293\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12288\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12288\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12299\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__12296\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12293\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__12288\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__12279\,
            I => \N__12276\
        );

    \I__2083\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12268\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12268\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12263\
        );

    \I__2080\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12263\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12268\,
            I => \N__12259\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__12263\,
            I => \N__12256\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12253\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__12259\,
            I => \N__12250\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__12256\,
            I => \Lab_UT.didp.un24_ce_3\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__12253\,
            I => \Lab_UT.didp.un24_ce_3\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__12250\,
            I => \Lab_UT.didp.un24_ce_3\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12240\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12240\,
            I => \N__12237\
        );

    \I__2070\ : Span4Mux_h
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__12234\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12228\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12228\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12222\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__12216\,
            I => \N__12213\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__12210\,
            I => \uu2.N_149\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__12204\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12195\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12195\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12189\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12189\,
            I => \uu2.N_25\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12177\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12177\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12177\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12177\,
            I => \Lab_UT.didp.countrce1.ce_12_1_1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12170\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12166\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12170\,
            I => \N__12163\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12160\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12166\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__12163\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12160\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__2039\ : Span4Mux_v
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__12141\,
            I => \Lab_UT.didp.countrce4.un20_qPone\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12132\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12132\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12128\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12124\
        );

    \I__2033\ : Span4Mux_s2_v
    port map (
            O => \N__12128\,
            I => \N__12121\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12118\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12124\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__12121\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12118\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12108\,
            I => \N__12103\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12100\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12096\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__12103\,
            I => \N__12088\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12100\,
            I => \N__12085\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__12099\,
            I => \N__12081\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12096\,
            I => \N__12076\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__12095\,
            I => \N__12073\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \N__12069\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \N__12066\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__12092\,
            I => \N__12063\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12060\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__12088\,
            I => \N__12057\
        );

    \I__2014\ : Span4Mux_s2_v
    port map (
            O => \N__12085\,
            I => \N__12054\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12045\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12045\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12045\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12045\
        );

    \I__2009\ : Span4Mux_s2_v
    port map (
            O => \N__12076\,
            I => \N__12042\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12033\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12033\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12033\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12033\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12028\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12028\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__12057\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__12054\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12045\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__12042\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12033\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12028\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12012\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12012\,
            I => \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__12009\,
            I => \N__12006\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12000\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12005\,
            I => \N__12000\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12000\,
            I => \N__11997\
        );

    \I__1990\ : Span4Mux_s2_v
    port map (
            O => \N__11997\,
            I => \N__11994\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__11994\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11988\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11988\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__11985\,
            I => \N__11982\
        );

    \I__1985\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11979\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11979\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11973\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__11973\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11970\,
            I => \N__11967\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__11967\,
            I => \N__11964\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__11964\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__11961\,
            I => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11955\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__11955\,
            I => \uu2.N_14\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11949\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11949\,
            I => \N__11946\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__11946\,
            I => \uu2.bitmap_RNI2Q8F1Z0Z_111\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11940\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__11940\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11930\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11927\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11920\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11920\
        );

    \I__1966\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11920\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__11930\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11927\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__11920\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11910\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11910\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1960\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11904\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__11904\,
            I => \uu2.N_166\
        );

    \I__1958\ : CEMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__11898\,
            I => \N__11894\
        );

    \I__1956\ : CEMux
    port map (
            O => \N__11897\,
            I => \N__11891\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__11894\,
            I => \N__11887\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__11891\,
            I => \N__11884\
        );

    \I__1953\ : CEMux
    port map (
            O => \N__11890\,
            I => \N__11881\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__11887\,
            I => \N__11878\
        );

    \I__1951\ : Span4Mux_s0_v
    port map (
            O => \N__11884\,
            I => \N__11875\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__11881\,
            I => \N__11872\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__11878\,
            I => \uu2.N_33_1\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__11875\,
            I => \uu2.N_33_1\
        );

    \I__1947\ : Odrv12
    port map (
            O => \N__11872\,
            I => \uu2.N_33_1\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11859\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__1943\ : Span4Mux_s0_v
    port map (
            O => \N__11856\,
            I => \N__11853\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__11853\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__11850\,
            I => \N__11847\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11844\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__11844\,
            I => \N__11841\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__11841\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__11838\,
            I => \N__11835\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11829\
        );

    \I__1934\ : Odrv12
    port map (
            O => \N__11829\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__11826\,
            I => \N__11823\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11820\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1930\ : Odrv12
    port map (
            O => \N__11817\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11811\,
            I => \Lab_UT.dictrl.g1_0Z0Z_5\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__11808\,
            I => \Lab_UT.dictrl.g1_0_4_0_cascade_\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11802\,
            I => \Lab_UT.dictrl.g0_5_4_0\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__11799\,
            I => \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__11796\,
            I => \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11790\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__11790\,
            I => \Lab_UT.dictrl.g0_5_3_0\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__11787\,
            I => \Lab_UT.dictrl.G_25_i_o3_3_cascade_\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11781\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__11781\,
            I => \Lab_UT.dictrl.alarmstate8Z0Z_3\
        );

    \I__1917\ : CEMux
    port map (
            O => \N__11778\,
            I => \N__11775\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__11772\,
            I => \Lab_UT.didp.regrce2.LdAStens_0\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__11769\,
            I => \N__11765\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__11768\,
            I => \N__11762\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11757\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11757\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__11754\,
            I => \N__11750\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11747\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__11750\,
            I => \Lab_UT.dictrl.alarmstateZ0Z8\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11747\,
            I => \Lab_UT.dictrl.alarmstateZ0Z8\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__11742\,
            I => \N__11739\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__11733\,
            I => \Lab_UT.dictrl.m37_N_2LZ0Z1\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__11730\,
            I => \Lab_UT.didp.countrce4.q_5_3_cascade_\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11724\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__11721\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_2\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11715\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_2_2\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \Lab_UT.didp.countrce4.q_5_0_cascade_\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__11709\,
            I => \N__11705\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__11708\,
            I => \N__11694\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11690\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11685\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11685\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11680\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11680\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11671\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11671\
        );

    \I__1885\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11671\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11697\,
            I => \N__11671\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11666\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11666\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__11690\,
            I => \G_181\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11685\,
            I => \G_181\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__11680\,
            I => \G_181\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11671\,
            I => \G_181\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11666\,
            I => \G_181\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11638\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11638\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11638\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11633\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11633\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11630\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11625\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11625\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11622\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11619\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11616\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11638\,
            I => \G_179\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11633\,
            I => \G_179\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__11630\,
            I => \G_179\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11625\,
            I => \G_179\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11622\,
            I => \G_179\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11619\,
            I => \G_179\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__11616\,
            I => \G_179\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__11601\,
            I => \N__11598\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11595\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__11595\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__11592\,
            I => \N__11588\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__11591\,
            I => \N__11584\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11574\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11574\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11574\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11571\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11568\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11565\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11562\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11571\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11568\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11565\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__11562\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__11553\,
            I => \N__11548\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11545\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11541\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11538\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__11545\,
            I => \N__11535\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11532\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11541\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__11538\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__11535\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11532\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \N__11520\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11517\,
            I => \Lab_UT.dispString.N_140\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__11514\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11508\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11508\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11502\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11502\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11490\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11483\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11483\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11483\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11478\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11478\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__11478\,
            I => \N__11475\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__11475\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__11472\,
            I => \N__11469\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11466\,
            I => \Lab_UT.didp.countrce1.un20_qPone\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \Lab_UT.didp.countrce1.q_5_3_cascade_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11457\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__1809\ : Span4Mux_h
    port map (
            O => \N__11454\,
            I => \N__11451\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__11451\,
            I => \Lab_UT.dispString.N_137\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11445\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11445\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11439\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11439\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11430\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11430\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__11430\,
            I => \N__11425\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11420\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11420\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__11425\,
            I => \Lab_UT.didp.ce_12_1\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__11420\,
            I => \Lab_UT.didp.ce_12_1\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \Lab_UT.didp.ce_12_1_cascade_\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \Lab_UT.didp.ce_12_3_cascade_\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11406\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11406\,
            I => \N__11403\
        );

    \I__1792\ : Span4Mux_h
    port map (
            O => \N__11403\,
            I => \N__11400\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__11400\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_1\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__11397\,
            I => \N__11389\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11385\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11382\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11371\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11371\
        );

    \I__1785\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11371\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11371\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11371\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11385\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__11382\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11371\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__11364\,
            I => \uu2.N_24_cascade_\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11358\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11358\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11349\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11349\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11342\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11339\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__11342\,
            I => \uu2.N_31_i\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11339\,
            I => \uu2.N_31_i\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__11334\,
            I => \uu2.N_26_cascade_\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11328\,
            I => \uu2.bitmap_pmux_27_ns_1\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11322\,
            I => \uu2.N_404\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11319\,
            I => \N__11315\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__11318\,
            I => \N__11312\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11306\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11306\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11303\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__11306\,
            I => \N__11298\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__11303\,
            I => \N__11298\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__11298\,
            I => \uu2.un51_w_data_displaying_i_a2_1\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__11295\,
            I => \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11292\,
            I => \N__11286\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11286\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__11286\,
            I => \N__11283\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__11283\,
            I => \uu2.w_data_displaying_2_i_a2_i_a3_2_0\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11276\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11273\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11276\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__11273\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11265\,
            I => \N__11262\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__11262\,
            I => \uu2.w_addr_displaying_RNI03P31Z0Z_4\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11259\,
            I => \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11253\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11250\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__11250\,
            I => \uu2.bitmap_pmux_sn_i7_mux_0\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11229\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11229\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11229\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11229\
        );

    \I__1736\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11229\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11229\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11229\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__1733\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11223\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11223\,
            I => \G_180\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11220\,
            I => \Lab_UT.dictrl.alarmstate_1_0_cascade_\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11210\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11210\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11207\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11210\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11207\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__11202\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11195\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11192\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11195\,
            I => \G_184\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__11192\,
            I => \G_184\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11187\,
            I => \resetGen.escKeyZ0Z_5_cascade_\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11178\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11178\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__11178\,
            I => \N__11172\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11165\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11165\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11165\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__11172\,
            I => \N__11160\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__11165\,
            I => \N__11160\
        );

    \I__1711\ : Span4Mux_h
    port map (
            O => \N__11160\,
            I => \N__11157\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__11157\,
            I => \resetGen.escKeyZ0\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11151\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11151\,
            I => \resetGen.escKeyZ0Z_4\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11143\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11140\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11137\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11143\,
            I => \N__11134\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11140\,
            I => \G_186\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11137\,
            I => \G_186\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__11134\,
            I => \G_186\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11124\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11120\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \N__11117\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__11120\,
            I => \N__11113\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11110\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11107\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__11113\,
            I => \L3_tx_data_6\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11110\,
            I => \L3_tx_data_6\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11107\,
            I => \L3_tx_data_6\
        );

    \I__1691\ : SRMux
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11091\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__11096\,
            I => \N__11088\
        );

    \I__1688\ : IoInMux
    port map (
            O => \N__11095\,
            I => \N__11085\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11082\
        );

    \I__1686\ : Span4Mux_s3_h
    port map (
            O => \N__11091\,
            I => \N__11079\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11076\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11073\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11082\,
            I => \N__11070\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__11079\,
            I => \N__11065\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11076\,
            I => \N__11065\
        );

    \I__1680\ : Span12Mux_s5_v
    port map (
            O => \N__11073\,
            I => \N__11062\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__11070\,
            I => \N__11059\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__11065\,
            I => \N__11056\
        );

    \I__1677\ : Odrv12
    port map (
            O => \N__11062\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__11059\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__11056\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11045\
        );

    \I__1673\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11042\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11045\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11042\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__11037\,
            I => \Lab_UT.un1_idle_4_0_iclkZ0_cascade_\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__11031\,
            I => \G_185\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__11028\,
            I => \G_185_cascade_\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__11025\,
            I => \Lab_UT.dispString.N_117_cascade_\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11019\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__1663\ : Span4Mux_s1_v
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__11013\,
            I => \N__11008\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11003\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11003\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__11008\,
            I => \L3_tx_data_1\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11003\,
            I => \L3_tx_data_1\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10995\,
            I => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__10992\,
            I => \G_180_cascade_\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__10989\,
            I => \G_181_cascade_\
        );

    \I__1653\ : CEMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10980\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__10977\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__10974\,
            I => \N__10971\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__10968\,
            I => \uu2.un1_w_user_lfZ0Z_4\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10961\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__10964\,
            I => \N__10958\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10954\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10949\
        );

    \I__1642\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10949\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__10954\,
            I => \L3_tx_data_5\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__10949\,
            I => \L3_tx_data_5\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__10944\,
            I => \N__10940\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10936\
        );

    \I__1637\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10931\
        );

    \I__1636\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10931\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__10936\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__10931\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10920\
        );

    \I__1631\ : Odrv12
    port map (
            O => \N__10920\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_3\
        );

    \I__1630\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10914\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__10914\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_3\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10908\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__10908\,
            I => \uu2.un1_w_user_lfZ0Z_3\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10902\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10899\
        );

    \I__1624\ : Span4Mux_s3_v
    port map (
            O => \N__10899\,
            I => \N__10894\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10889\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10889\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__10894\,
            I => \L3_tx_data_3\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__10889\,
            I => \L3_tx_data_3\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10881\,
            I => \N__10878\
        );

    \I__1617\ : Span4Mux_s3_v
    port map (
            O => \N__10878\,
            I => \N__10873\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10868\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10868\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__10873\,
            I => \L3_tx_data_0\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10868\,
            I => \L3_tx_data_0\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10858\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10853\
        );

    \I__1610\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10853\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__10858\,
            I => \uu2.un1_w_user_crZ0Z_3\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10853\,
            I => \uu2.un1_w_user_crZ0Z_3\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10845\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10845\,
            I => \Lab_UT.dispString.dOutP_1_iv_i_1_4\
        );

    \I__1605\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10839\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10836\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__10836\,
            I => \N__10831\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10826\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10826\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__10831\,
            I => \L3_tx_data_4\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10826\,
            I => \L3_tx_data_4\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10815\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10815\,
            I => \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__10812\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10803\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__10803\,
            I => \N__10800\
        );

    \I__1591\ : Odrv12
    port map (
            O => \N__10800\,
            I => \uu2.un20_w_addr_userZ0Z_1\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10793\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10789\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__10793\,
            I => \N__10786\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10783\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10789\,
            I => \L3_tx_data_rdy\
        );

    \I__1585\ : Odrv12
    port map (
            O => \N__10786\,
            I => \L3_tx_data_rdy\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10783\,
            I => \L3_tx_data_rdy\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__10776\,
            I => \Lab_UT.dispString.N_124_cascade_\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__10773\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10767\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__10767\,
            I => \uu2.bitmap_pmux_sn_i5_mux\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10761\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__10761\,
            I => \uu2.bitmap_pmux_u_1\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10754\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10751\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__10754\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10751\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1573\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10743\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10743\,
            I => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10737\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__10737\,
            I => \uu2.w_addr_displaying_RNI0NG56Z0Z_4\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10730\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10727\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10724\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__10727\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__10724\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__1562\ : Odrv12
    port map (
            O => \N__10713\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10707\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__10707\,
            I => \uu2.N_401\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__10704\,
            I => \uu2.N_406_cascade_\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10695\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__10695\,
            I => \uu2.bitmap_pmux\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__10692\,
            I => \uu2.N_383_cascade_\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__10689\,
            I => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10683\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__10683\,
            I => \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\
        );

    \I__1551\ : CEMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10674\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__10674\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__10671\,
            I => \uu2.un28_w_addr_user_i_cascade_\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__10668\,
            I => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__10665\,
            I => \uu2.bitmap_pmux_sn_N_15_cascade_\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__10662\,
            I => \G_182_cascade_\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10654\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10649\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10649\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10654\,
            I => \G_187\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__10649\,
            I => \G_187\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__10644\,
            I => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10632\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10632\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10632\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10632\,
            I => \G_183\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10623\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10623\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__10623\,
            I => \G_182\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10611\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10611\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10618\,
            I => \N__10606\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10606\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10603\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10611\,
            I => \N__10600\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10596\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10603\,
            I => \N__10593\
        );

    \I__1523\ : Span4Mux_s3_h
    port map (
            O => \N__10600\,
            I => \N__10590\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10587\
        );

    \I__1521\ : Span12Mux_s5_v
    port map (
            O => \N__10596\,
            I => \N__10582\
        );

    \I__1520\ : Span12Mux_s3_h
    port map (
            O => \N__10593\,
            I => \N__10582\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__10590\,
            I => \N__10579\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__10587\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1517\ : Odrv12
    port map (
            O => \N__10582\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__10579\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10569\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10566\
        );

    \I__1513\ : Span4Mux_h
    port map (
            O => \N__10566\,
            I => \N__10563\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__10563\,
            I => vbuf_tx_data_6
        );

    \I__1511\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10551\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__10551\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10545\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10542\
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__10542\,
            I => vbuf_tx_data_7
        );

    \I__1504\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__10536\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__10533\,
            I => \N__10530\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10527\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10524\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__10524\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__1498\ : SRMux
    port map (
            O => \N__10521\,
            I => \N__10518\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10514\
        );

    \I__1496\ : CEMux
    port map (
            O => \N__10517\,
            I => \N__10511\
        );

    \I__1495\ : Span4Mux_s3_v
    port map (
            O => \N__10514\,
            I => \N__10508\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10511\,
            I => \N__10505\
        );

    \I__1493\ : Span4Mux_h
    port map (
            O => \N__10508\,
            I => \N__10500\
        );

    \I__1492\ : Span4Mux_s3_v
    port map (
            O => \N__10505\,
            I => \N__10500\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__10500\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10494\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10494\,
            I => \G_188\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__10491\,
            I => \G_188_cascade_\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10485\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__10485\,
            I => \Lab_UT.un1_rst_0_iclkZ0\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__10482\,
            I => \N__10479\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10473\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10468\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10468\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__10476\,
            I => \N__10465\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10462\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10468\,
            I => \N__10459\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10456\
        );

    \I__1477\ : Span4Mux_s3_h
    port map (
            O => \N__10462\,
            I => \N__10451\
        );

    \I__1476\ : Span4Mux_s1_v
    port map (
            O => \N__10459\,
            I => \N__10451\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10456\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__10451\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10436\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10433\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10426\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10426\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10426\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__10436\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10433\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10426\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10419\,
            I => \N__10416\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10412\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__10415\,
            I => \N__10409\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10406\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10403\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__10406\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10403\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10395\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10395\,
            I => \N__10392\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__10392\,
            I => \N__10385\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10376\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10376\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10376\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10376\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__10385\,
            I => \uu2.un306_ci\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10376\,
            I => \uu2.un306_ci\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10367\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10364\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10360\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10357\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10354\
        );

    \I__1443\ : Span4Mux_s2_h
    port map (
            O => \N__10360\,
            I => \N__10349\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10349\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__10354\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__10349\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10338\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10338\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10338\,
            I => \N__10335\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__10332\,
            I => \uu2.un284_ci\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__10329\,
            I => \N__10324\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10320\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10315\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10315\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__10323\,
            I => \N__10312\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10306\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10306\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10301\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10301\
        );

    \I__1425\ : Span4Mux_s3_h
    port map (
            O => \N__10306\,
            I => \N__10298\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10301\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__10298\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10287\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10287\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10287\,
            I => \uu2.N_31\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10284\,
            I => \uu2.N_31_cascade_\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10278\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10278\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__10275\,
            I => \N__10270\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10264\
        );

    \I__1414\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10264\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10261\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10258\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10255\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__10261\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10258\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__10255\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__10248\,
            I => \N__10244\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \N__10239\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10235\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10230\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10230\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10225\
        );

    \I__1401\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10225\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10220\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10220\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10225\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__10220\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__10215\,
            I => \N__10210\
        );

    \I__1395\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10202\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10202\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10199\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10192\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10192\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10192\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10202\,
            I => \N__10189\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10199\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10192\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__10189\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1385\ : CEMux
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10179\,
            I => \N__10176\
        );

    \I__1383\ : Span4Mux_s1_v
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__10173\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10164\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10161\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10156\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10156\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10164\,
            I => \N__10153\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__10161\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10156\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__10153\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10135\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10124\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10124\
        );

    \I__1369\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10124\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10124\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10124\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__10135\,
            I => \N__10119\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10119\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__10119\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10107\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10101\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10101\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10098\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10107\,
            I => \N__10095\
        );

    \I__1357\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10092\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10101\,
            I => \N__10089\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__10098\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__10095\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__10092\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__10089\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10077\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10073\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10070\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__10073\,
            I => \N__10063\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10070\,
            I => \N__10063\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10058\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10058\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__10063\,
            I => \uu2.un404_ci_0\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__10058\,
            I => \uu2.un404_ci_0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__10053\,
            I => \uu2.un404_ci_0_cascade_\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__10050\,
            I => \N__10047\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10042\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10039\
        );

    \I__1338\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10036\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__10042\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10039\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__10036\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__10029\,
            I => \N__10025\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__10028\,
            I => \N__10021\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10017\
        );

    \I__1331\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10010\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10010\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10010\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10017\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__10010\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10005\,
            I => \N__10002\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10002\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9996\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__9996\,
            I => \uu2.mem0.w_data_6\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__9990\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9984\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__9984\,
            I => \uu2.N_34\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__9981\,
            I => \uu2.N_34_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9975\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__9975\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9969\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__9969\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9963\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9963\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9955\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9952\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9949\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__9955\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__9952\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__9949\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1305\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__9939\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9936\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9929\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9926\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9929\,
            I => \N__9923\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9926\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__9923\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9918\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__9915\,
            I => \N__9912\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9907\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9904\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9901\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9907\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9904\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__9901\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9891\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9888\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9879\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9872\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9872\
        );

    \I__1283\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9872\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__9879\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__9872\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__9867\,
            I => \N__9861\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9855\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9852\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9849\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9841\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9838\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9833\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9833\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9826\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9826\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9826\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9815\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9815\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9815\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9815\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9815\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9841\,
            I => \buart.Z_rx.startbit\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__9838\,
            I => \buart.Z_rx.startbit\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__9833\,
            I => \buart.Z_rx.startbit\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__9826\,
            I => \buart.Z_rx.startbit\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9815\,
            I => \buart.Z_rx.startbit\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9804\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__9801\,
            I => \N__9797\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__9800\,
            I => \N__9794\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9791\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9788\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9791\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9788\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__9783\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9773\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9770\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9773\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__9770\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9762\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9762\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__9759\,
            I => \N__9754\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__9758\,
            I => \N__9751\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__9757\,
            I => \N__9748\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9745\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9740\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9740\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9745\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9740\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9732\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__9729\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9720\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9716\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9711\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9711\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__9720\,
            I => \N__9708\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9705\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9716\,
            I => \N__9700\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9711\,
            I => \N__9700\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__9708\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__9705\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__9700\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1222\ : IoInMux
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__1220\ : Span4Mux_s2_v
    port map (
            O => \N__9687\,
            I => \N__9684\
        );

    \I__1219\ : Span4Mux_h
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__9681\,
            I => \buart.Z_rx.sample\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__9678\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__9675\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9664\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9659\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9659\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__9664\,
            I => \buart.Z_rx.idle\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9659\,
            I => \buart.Z_rx.idle\
        );

    \I__1209\ : CEMux
    port map (
            O => \N__9654\,
            I => \N__9648\
        );

    \I__1208\ : CEMux
    port map (
            O => \N__9653\,
            I => \N__9645\
        );

    \I__1207\ : CEMux
    port map (
            O => \N__9652\,
            I => \N__9642\
        );

    \I__1206\ : CEMux
    port map (
            O => \N__9651\,
            I => \N__9639\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9648\,
            I => \N__9634\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__9645\,
            I => \N__9634\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9631\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9628\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__9634\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1200\ : Odrv12
    port map (
            O => \N__9631\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__9628\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9616\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9611\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9611\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9616\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__9611\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__9606\,
            I => \N__9602\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9605\,
            I => \N__9599\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9594\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9587\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9587\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9587\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9594\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9587\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__9582\,
            I => \N__9579\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9576\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9576\,
            I => \N__9573\
        );

    \I__1182\ : Span12Mux_s9_v
    port map (
            O => \N__9573\,
            I => \N__9570\
        );

    \I__1181\ : Odrv12
    port map (
            O => \N__9570\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9563\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9552\
        );

    \I__1176\ : Span4Mux_v
    port map (
            O => \N__9557\,
            I => \N__9552\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__9552\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9542\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__9545\,
            I => \N__9537\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9533\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9530\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9527\
        );

    \I__1168\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9522\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9522\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__9533\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9530\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__9527\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9522\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__9513\,
            I => \resetGen.un241_ci_cascade_\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9505\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9500\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9500\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__9505\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9500\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__9495\,
            I => \N__9492\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9484\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9484\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9479\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9479\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9484\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9479\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__9474\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9465\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9465\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9465\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1145\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9453\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9453\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9453\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9453\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9447\,
            I => \resetGen.un241_ci\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__9444\,
            I => \resetGen.reset_count_2_0_4_cascade_\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9431\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9431\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9424\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9424\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9424\
        );

    \I__1133\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9421\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9431\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9424\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__9421\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9410\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9407\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9410\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__9407\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9394\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9391\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9388\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9394\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9391\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__9388\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__9381\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9368\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9368\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9368\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9365\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9368\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9365\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9357\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9357\,
            I => \uu0.un4_l_count_16\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9347\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9340\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9340\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9340\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9336\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9347\,
            I => \N__9331\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9331\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9328\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9325\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__9331\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9328\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__9325\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__9318\,
            I => \N__9314\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9308\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9301\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9301\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9301\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9298\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9308\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9301\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__9298\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__9291\,
            I => \CONSTANT_ONE_NET_cascade_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9285\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9285\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9272\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9272\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9272\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9269\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9272\,
            I => \N__9265\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9262\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9259\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__9265\,
            I => \N__9256\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__9262\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__9259\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__9256\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__9243\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9236\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9233\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9230\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__9233\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__9230\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9210\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9203\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9203\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9203\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9200\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9197\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9192\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9192\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9189\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9186\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9183\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9178\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9178\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9210\,
            I => \N__9175\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9203\,
            I => \uu0.un4_l_count_0\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__9200\,
            I => \uu0.un4_l_count_0\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9197\,
            I => \uu0.un4_l_count_0\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9192\,
            I => \uu0.un4_l_count_0\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__9189\,
            I => \uu0.un4_l_count_0\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9186\,
            I => \uu0.un4_l_count_0\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__9183\,
            I => \uu0.un4_l_count_0\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9178\,
            I => \uu0.un4_l_count_0\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9175\,
            I => \uu0.un4_l_count_0\
        );

    \I__1043\ : IoInMux
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__1041\ : Span4Mux_s1_h
    port map (
            O => \N__9150\,
            I => \N__9147\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__9147\,
            I => \uu0.un11_l_count_i\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__9144\,
            I => \uu0.un143_ci_0_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__9141\,
            I => \N__9131\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__9140\,
            I => \N__9128\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__9139\,
            I => \N__9125\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9118\
        );

    \I__1034\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9118\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9109\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9109\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9109\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9109\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9100\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9100\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9100\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9100\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9118\,
            I => \uu0.un110_ci\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9109\,
            I => \uu0.un110_ci\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9100\,
            I => \uu0.un110_ci\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9085\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9074\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9074\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9074\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9074\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9074\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9085\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9074\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1014\ : CEMux
    port map (
            O => \N__9069\,
            I => \N__9057\
        );

    \I__1013\ : CEMux
    port map (
            O => \N__9068\,
            I => \N__9057\
        );

    \I__1012\ : CEMux
    port map (
            O => \N__9067\,
            I => \N__9057\
        );

    \I__1011\ : CEMux
    port map (
            O => \N__9066\,
            I => \N__9057\
        );

    \I__1010\ : GlobalMux
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__1009\ : gio2CtrlBuf
    port map (
            O => \N__9054\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__9051\,
            I => \N__9046\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__9050\,
            I => \N__9042\
        );

    \I__1006\ : InMux
    port map (
            O => \N__9049\,
            I => \N__9039\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9032\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9032\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9032\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9029\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9032\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__9029\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__9024\,
            I => \N__9020\
        );

    \I__998\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9016\
        );

    \I__997\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9013\
        );

    \I__996\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9010\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9016\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__9013\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9010\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8996\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__9002\,
            I => \N__8993\
        );

    \I__990\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8984\
        );

    \I__989\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8984\
        );

    \I__988\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8984\
        );

    \I__987\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8984\
        );

    \I__986\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8981\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__8984\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__8981\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__983\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8973\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8973\,
            I => \uu0.un4_l_count_12\
        );

    \I__981\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8967\,
            I => \uu0.un4_l_count_18\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__8964\,
            I => \uu0.un4_l_count_13_cascade_\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__8961\,
            I => \N__8957\
        );

    \I__977\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8946\
        );

    \I__976\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8946\
        );

    \I__975\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8946\
        );

    \I__974\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8946\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__8946\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__972\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8936\
        );

    \I__971\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8936\
        );

    \I__970\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8933\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8936\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8933\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__8928\,
            I => \N__8923\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__8927\,
            I => \N__8920\
        );

    \I__965\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8913\
        );

    \I__964\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8913\
        );

    \I__963\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8913\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__8913\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__961\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8900\
        );

    \I__960\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8900\
        );

    \I__959\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8900\
        );

    \I__958\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8897\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__8900\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8897\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__955\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8889\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8889\,
            I => \uu0.un187_ci_1\
        );

    \I__953\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8877\
        );

    \I__952\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8877\
        );

    \I__951\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8877\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__8877\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__949\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8863\
        );

    \I__948\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8863\
        );

    \I__947\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8863\
        );

    \I__946\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8858\
        );

    \I__945\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8858\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8855\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__8858\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__8855\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__940\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8841\
        );

    \I__939\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8838\
        );

    \I__938\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8833\
        );

    \I__937\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8833\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8828\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8828\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__8833\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__8828\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__8823\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__8820\,
            I => \N__8816\
        );

    \I__930\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8811\
        );

    \I__929\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8804\
        );

    \I__928\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8804\
        );

    \I__927\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8804\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8801\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8804\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__8801\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__922\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8787\
        );

    \I__921\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8784\
        );

    \I__920\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8779\
        );

    \I__919\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8779\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8787\,
            I => \uu0.un154_ci_9\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__8784\,
            I => \uu0.un154_ci_9\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__8779\,
            I => \uu0.un154_ci_9\
        );

    \I__915\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8764\
        );

    \I__914\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8764\
        );

    \I__913\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8759\
        );

    \I__912\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8759\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8764\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8759\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__8754\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__8751\,
            I => \N__8745\
        );

    \I__907\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8742\
        );

    \I__906\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8739\
        );

    \I__905\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8736\
        );

    \I__904\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8733\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8742\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8739\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8736\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8733\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__898\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8710\
        );

    \I__897\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8710\
        );

    \I__896\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8710\
        );

    \I__895\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8705\
        );

    \I__894\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8705\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8710\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8705\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__891\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8688\
        );

    \I__890\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8688\
        );

    \I__889\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8688\
        );

    \I__888\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8688\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8688\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \uu2.vbuf_count.un328_ci_3_cascade_\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__8682\,
            I => \N__8677\
        );

    \I__884\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8674\
        );

    \I__883\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8669\
        );

    \I__882\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8669\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8674\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8669\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__8664\,
            I => \N__8658\
        );

    \I__878\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8646\
        );

    \I__877\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8646\
        );

    \I__876\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8646\
        );

    \I__875\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8646\
        );

    \I__874\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8646\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8646\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__872\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8636\
        );

    \I__871\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8636\
        );

    \I__870\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8633\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8636\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__8633\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__866\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8620\
        );

    \I__865\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8617\
        );

    \I__864\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8614\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8620\,
            I => \N__8611\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8617\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8614\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__8611\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__8604\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8598\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__856\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8591\
        );

    \I__855\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8588\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8585\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__8588\,
            I => \N__8582\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__8585\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__8582\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__850\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8568\
        );

    \I__849\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8568\
        );

    \I__848\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8568\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__8565\,
            I => \uu0.un198_ci_2\
        );

    \I__845\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8559\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__842\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8550\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__840\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8542\
        );

    \I__839\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8537\
        );

    \I__838\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8537\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8542\,
            I => \N__8534\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8537\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__8534\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__8529\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__833\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8522\
        );

    \I__832\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8519\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8522\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8519\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__829\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8511\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__827\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8505\,
            I => \uu2.un350_ci\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8502\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__824\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8496\,
            I => vbuf_tx_data_0
        );

    \I__822\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8490\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__820\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8484\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__816\ : Span12Mux_s1_h
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__8472\,
            I => o_serial_data_c
        );

    \I__814\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8466\,
            I => vbuf_tx_data_1
        );

    \I__812\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8460\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8460\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__810\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8454\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8454\,
            I => vbuf_tx_data_2
        );

    \I__808\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8448\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__806\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8442\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8442\,
            I => vbuf_tx_data_3
        );

    \I__804\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8436\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__802\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8430\,
            I => vbuf_tx_data_4
        );

    \I__800\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8424\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__798\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8418\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8418\,
            I => vbuf_tx_data_5
        );

    \I__796\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8412\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8412\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__794\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8403\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__8403\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__791\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8396\
        );

    \I__790\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8390\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8396\,
            I => \N__8387\
        );

    \I__788\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8380\
        );

    \I__787\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8380\
        );

    \I__786\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8380\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8390\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__8387\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8380\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__782\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8370\,
            I => \uu2.r_data_wire_0\
        );

    \I__780\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__8364\,
            I => \uu2.r_data_wire_1\
        );

    \I__778\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8358\,
            I => \uu2.r_data_wire_2\
        );

    \I__776\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8352\,
            I => \uu2.r_data_wire_3\
        );

    \I__774\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8346\,
            I => \uu2.r_data_wire_4\
        );

    \I__772\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8340\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8340\,
            I => \uu2.r_data_wire_5\
        );

    \I__770\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8334\,
            I => \uu2.r_data_wire_6\
        );

    \I__768\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__8328\,
            I => \uu2.r_data_wire_7\
        );

    \I__766\ : InMux
    port map (
            O => \N__8325\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__765\ : InMux
    port map (
            O => \N__8322\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__764\ : InMux
    port map (
            O => \N__8319\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__8316\,
            I => \buart.Z_rx.valid_0_cascade_\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__761\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8304\
        );

    \I__760\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8297\
        );

    \I__759\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8297\
        );

    \I__758\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8297\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8304\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__8297\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__8292\,
            I => \buart.Z_rx.idle_0_cascade_\
        );

    \I__754\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8286\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__8283\,
            I => \N__8278\
        );

    \I__751\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8273\
        );

    \I__750\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8264\
        );

    \I__749\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8264\
        );

    \I__748\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8264\
        );

    \I__747\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8264\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8273\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8264\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__8259\,
            I => \N__8254\
        );

    \I__743\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8251\
        );

    \I__742\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8248\
        );

    \I__741\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8245\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8251\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8248\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8245\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__8235\,
            I => \N__8231\
        );

    \I__735\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8226\
        );

    \I__734\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8221\
        );

    \I__733\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8221\
        );

    \I__732\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8218\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8213\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8221\,
            I => \N__8213\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8218\,
            I => \uu0.un66_ci\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__8213\,
            I => \uu0.un66_ci\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__8208\,
            I => \N__8203\
        );

    \I__726\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8196\
        );

    \I__725\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8196\
        );

    \I__724\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8196\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8196\,
            I => \N__8193\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__8193\,
            I => \uu0.un88_ci_3\
        );

    \I__721\ : InMux
    port map (
            O => \N__8190\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__720\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8178\
        );

    \I__719\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8178\
        );

    \I__718\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8178\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8178\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__8175\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__714\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8166\,
            I => \uu0.un99_ci_0\
        );

    \I__712\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8158\
        );

    \I__711\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8153\
        );

    \I__710\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8153\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8158\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__8153\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__707\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8145\,
            I => \uu0.un44_ci\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__8142\,
            I => \uu0.un44_ci_cascade_\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__8139\,
            I => \uu0.un165_ci_0_cascade_\
        );

    \I__703\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8130\
        );

    \I__702\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8130\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__8130\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__8127\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__699\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8115\
        );

    \I__698\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8115\
        );

    \I__697\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8115\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8115\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__695\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__693\ : IoSpan4Mux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__692\ : IoSpan4Mux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__8100\,
            I => \uart_RXD\
        );

    \I__690\ : IoInMux
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__688\ : Span12Mux_s5_v
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__687\ : Odrv12
    port map (
            O => \N__8088\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__686\ : IoInMux
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__684\ : IoSpan4Mux
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__8076\,
            I => clk_in_c
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__22262\
        );

    \INVuu2.w_addr_displaying_7C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_7C_net\,
            I => \N__22266\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__22270\
        );

    \INVuu2.bitmap_215C\ : INV
    port map (
            O => \INVuu2.bitmap_215C_net\,
            I => \N__22248\
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__22261\
        );

    \INVuu2.w_addr_displaying_fast_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_8C_net\,
            I => \N__22265\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__22240\
        );

    \INVuu2.bitmap_197C\ : INV
    port map (
            O => \INVuu2.bitmap_197C_net\,
            I => \N__22247\
        );

    \INVuu2.bitmap_168C\ : INV
    port map (
            O => \INVuu2.bitmap_168C_net\,
            I => \N__22255\
        );

    \INVuu2.w_addr_displaying_ness_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_ness_6C_net\,
            I => \N__22260\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__22235\
        );

    \INVuu2.w_addr_displaying_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_3C_net\,
            I => \N__22243\
        );

    \INVuu2.w_addr_user_2C\ : INV
    port map (
            O => \INVuu2.w_addr_user_2C_net\,
            I => \N__22250\
        );

    \INVuu2.vram_rd_clk_det_1C\ : INV
    port map (
            O => \INVuu2.vram_rd_clk_det_1C_net\,
            I => \N__22239\
        );

    \INVuu2.w_addr_displaying_1_rep1_nesrC\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            I => \N__22254\
        );

    \INVuu2.vram_rd_clk_det_0C\ : INV
    port map (
            O => \INVuu2.vram_rd_clk_det_0C_net\,
            I => \N__22246\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__22272\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8097\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9693\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9156\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14914\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8112\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22251\,
            ce => 'H',
            sr => \N__20679\
        );

    \uu0.l_count_RNIFAQ9_13_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8135\,
            in2 => \_gnd_net_\,
            in3 => \N__8122\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8206\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8794\,
            in2 => \_gnd_net_\,
            in3 => \N__8123\,
            lcout => OPEN,
            ltout => \uu0.un165_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_13_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8136\,
            in1 => \N__9137\,
            in2 => \N__8139\,
            in3 => \N__9223\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__9068\,
            sr => \N__20677\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8230\,
            in1 => \N__9376\,
            in2 => \N__8208\,
            in3 => \N__8163\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_12_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8124\,
            in1 => \N__8795\,
            in2 => \N__8127\,
            in3 => \N__9222\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__9068\,
            sr => \N__20677\
        );

    \uu0.l_count_6_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8207\,
            in1 => \N__9216\,
            in2 => \N__8235\,
            in3 => \N__9378\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__9068\,
            sr => \N__20677\
        );

    \uu0.l_count_15_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__8892\,
            in1 => \N__9138\,
            in2 => \N__9402\,
            in3 => \N__9224\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__9068\,
            sr => \N__20677\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8717\,
            in1 => \N__8161\,
            in2 => \N__8259\,
            in3 => \N__8185\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__9214\,
            in1 => \N__9124\,
            in2 => \N__9051\,
            in3 => \N__8576\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.l_count_17_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8577\,
            in1 => \N__9045\,
            in2 => \N__9139\,
            in3 => \N__8187\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8186\,
            in1 => \N__9123\,
            in2 => \N__9050\,
            in3 => \N__8575\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9213\,
            in2 => \N__8175\,
            in3 => \N__9414\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.l_count_3_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8258\,
            in1 => \N__8148\,
            in2 => \N__8850\,
            in3 => \N__9219\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.l_count_9_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__8718\,
            in1 => \_gnd_net_\,
            in2 => \N__9140\,
            in3 => \N__9093\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.l_count_7_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8162\,
            in1 => \N__8234\,
            in2 => \N__8172\,
            in3 => \N__9218\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22236\,
            ce => \N__9067\,
            sr => \N__20675\
        );

    \uu0.l_count_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9221\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => \N__9066\,
            sr => \N__20678\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__8909\,
            in1 => \N__8999\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.un44_ci\,
            ltout => \uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8142\,
            in3 => \N__8845\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => \N__9066\,
            sr => \N__20678\
        );

    \uu0.l_count_1_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__8910\,
            in1 => \N__9001\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => \N__9066\,
            sr => \N__20678\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8257\,
            in1 => \N__8844\,
            in2 => \N__9003\,
            in3 => \N__8908\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_4_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9215\,
            in2 => \N__8238\,
            in3 => \N__8815\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => \N__9066\,
            sr => \N__20678\
        );

    \uu0.l_count_5_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__8943\,
            in1 => \_gnd_net_\,
            in2 => \N__8820\,
            in3 => \N__8229\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => \N__9066\,
            sr => \N__20678\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8814\,
            in2 => \_gnd_net_\,
            in3 => \N__8942\,
            lcout => \uu0.un88_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__11184\,
            in1 => \N__9441\,
            in2 => \N__9495\,
            in3 => \N__9510\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__9440\,
            in1 => \N__9491\,
            in2 => \_gnd_net_\,
            in3 => \N__11183\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9436\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9719\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8400\,
            in2 => \_gnd_net_\,
            in3 => \N__8190\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9268\,
            in2 => \_gnd_net_\,
            in3 => \N__8325\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8282\,
            in2 => \_gnd_net_\,
            in3 => \N__8322\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__9540\,
            in1 => \N__9860\,
            in2 => \N__8313\,
            in3 => \N__8319\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22216\,
            ce => \N__9653\,
            sr => \N__20682\
        );

    \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8308\,
            in1 => \N__9281\,
            in2 => \N__8283\,
            in3 => \N__8394\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8307\,
            in2 => \_gnd_net_\,
            in3 => \N__9723\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8277\,
            in1 => \N__9280\,
            in2 => \N__8316\,
            in3 => \N__8393\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8276\,
            in2 => \_gnd_net_\,
            in3 => \N__8309\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9724\,
            in1 => \N__9282\,
            in2 => \N__8292\,
            in3 => \N__8395\,
            lcout => \buart.Z_rx.idle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001110100101110"
        )
    port map (
            in0 => \N__8281\,
            in1 => \N__9541\,
            in2 => \N__9867\,
            in3 => \N__8289\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22209\,
            ce => \N__9651\,
            sr => \N__20685\
        );

    \buart.Z_rx.bitcount_es_1_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__9864\,
            in1 => \N__8409\,
            in2 => \N__9549\,
            in3 => \N__8399\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22202\,
            ce => \N__9654\,
            sr => \N__20687\
        );

    \uu2.r_data_reg_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8349\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8343\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8337\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8331\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10680\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20418\,
            in1 => \N__8463\,
            in2 => \_gnd_net_\,
            in3 => \N__8499\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_0_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8493\,
            in2 => \_gnd_net_\,
            in3 => \N__20424\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.uart_tx_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8487\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_2_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8451\,
            in1 => \N__20421\,
            in2 => \_gnd_net_\,
            in3 => \N__8469\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_3_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20419\,
            in1 => \N__8439\,
            in2 => \_gnd_net_\,
            in3 => \N__8457\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_4_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__20422\,
            in2 => \_gnd_net_\,
            in3 => \N__8445\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_5_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20420\,
            in1 => \N__8415\,
            in2 => \_gnd_net_\,
            in3 => \N__8433\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \buart.Z_tx.shifter_6_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10560\,
            in1 => \N__20423\,
            in2 => \_gnd_net_\,
            in3 => \N__8421\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__20376\,
            sr => \N__20689\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8514\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__10169\,
            in1 => \N__8595\,
            in2 => \N__20438\,
            in3 => \N__20763\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8623\,
            in2 => \_gnd_net_\,
            in3 => \N__8508\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22258\,
            ce => 'H',
            sr => \N__20658\
        );

    \uu2.vram_rd_clk_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8547\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22258\,
            ce => 'H',
            sr => \N__20658\
        );

    \uu2.trig_rd_det_0_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10167\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22258\,
            ce => 'H',
            sr => \N__20658\
        );

    \uu2.trig_rd_det_1_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8526\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22258\,
            ce => 'H',
            sr => \N__20658\
        );

    \uu0.l_precount_0_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9339\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22258\,
            ce => 'H',
            sr => \N__20658\
        );

    \uu2.l_count_5_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10391\,
            in1 => \N__8663\,
            in2 => \_gnd_net_\,
            in3 => \N__8643\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \N__20686\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10442\,
            in1 => \N__10371\,
            in2 => \N__10415\,
            in3 => \N__10388\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__8546\,
            in1 => \N__8624\,
            in2 => \N__8502\,
            in3 => \N__8681\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \N__20686\
        );

    \uu2.l_count_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8662\,
            in1 => \N__10390\,
            in2 => \_gnd_net_\,
            in3 => \N__8545\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \N__20686\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8661\,
            in2 => \_gnd_net_\,
            in3 => \N__8642\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => \uu2.vbuf_count.un328_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_6_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10441\,
            in2 => \N__8685\,
            in3 => \N__10389\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \N__20686\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10439\,
            in1 => \N__8657\,
            in2 => \N__8682\,
            in3 => \N__10619\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_9_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10620\,
            in1 => \N__8680\,
            in2 => \N__8664\,
            in3 => \N__10440\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIFGGK1_3_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10370\,
            in1 => \N__8641\,
            in2 => \N__8628\,
            in3 => \N__8884\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10328\,
            in1 => \N__8873\,
            in2 => \N__8604\,
            in3 => \N__8601\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9398\,
            in1 => \N__8748\,
            in2 => \N__8796\,
            in3 => \N__8771\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8870\,
            in1 => \N__8562\,
            in2 => \N__8556\,
            in3 => \N__10327\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__10344\,
            in1 => \N__8871\,
            in2 => \N__8529\,
            in3 => \N__8886\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22245\,
            ce => 'H',
            sr => \N__20684\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8772\,
            in1 => \N__8793\,
            in2 => \_gnd_net_\,
            in3 => \N__8749\,
            lcout => \uu0.un187_ci_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8872\,
            in1 => \N__10616\,
            in2 => \N__10329\,
            in3 => \N__8885\,
            lcout => \uu2.un306_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10343\,
            in2 => \_gnd_net_\,
            in3 => \N__8874\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22245\,
            ce => 'H',
            sr => \N__20684\
        );

    \uu0.l_count_RNI04591_10_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8697\,
            in1 => \N__9088\,
            in2 => \N__8751\,
            in3 => \N__8846\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2GS72_4_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9350\,
            in1 => \N__8769\,
            in2 => \N__8823\,
            in3 => \N__8819\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_10_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8700\,
            in1 => \N__9092\,
            in2 => \N__8724\,
            in3 => \N__9136\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22237\,
            ce => \N__9069\,
            sr => \N__20680\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9089\,
            in1 => \N__8719\,
            in2 => \N__9024\,
            in3 => \N__8698\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8770\,
            in1 => \N__8750\,
            in2 => \N__8754\,
            in3 => \N__9135\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22237\,
            ce => \N__9069\,
            sr => \N__20680\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9090\,
            in1 => \N__8720\,
            in2 => \_gnd_net_\,
            in3 => \N__8699\,
            lcout => OPEN,
            ltout => \uu0.un143_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_11_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9023\,
            in1 => \N__9134\,
            in2 => \N__9144\,
            in3 => \N__9217\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22237\,
            ce => \N__9069\,
            sr => \N__20680\
        );

    \uu0.l_count_8_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__9091\,
            in1 => \_gnd_net_\,
            in2 => \N__9141\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22237\,
            ce => \N__9069\,
            sr => \N__20680\
        );

    \uu0.delay_line_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8956\,
            in1 => \N__9312\,
            in2 => \N__8928\,
            in3 => \N__9351\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => 'H',
            sr => \N__20676\
        );

    \uu0.l_count_RNI2CNU_11_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9049\,
            in1 => \N__9019\,
            in2 => \N__9002\,
            in3 => \N__8955\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_11_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8976\,
            in1 => \N__8970\,
            in2 => \N__8964\,
            in3 => \N__9360\,
            lcout => \uu0.un4_l_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_2_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9313\,
            in2 => \N__8961\,
            in3 => \N__9352\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => 'H',
            sr => \N__20676\
        );

    \uu0.l_precount_3_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9353\,
            in1 => \N__8926\,
            in2 => \N__9318\,
            in3 => \N__8960\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => 'H',
            sr => \N__20676\
        );

    \uu0.l_precount_RNI85Q91_3_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9311\,
            in1 => \N__8941\,
            in2 => \N__8927\,
            in3 => \N__8907\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI96A32_18_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9413\,
            in1 => \N__9397\,
            in2 => \N__9381\,
            in3 => \N__9375\,
            lcout => \uu0.un4_l_count_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22225\,
            ce => 'H',
            sr => \N__20681\
        );

    \buart.Z_rx.hh_1_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9566\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22225\,
            ce => 'H',
            sr => \N__20681\
        );

    \uu0.l_precount_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9354\,
            in2 => \_gnd_net_\,
            in3 => \N__9317\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22225\,
            ce => 'H',
            sr => \N__20681\
        );

    \uu0.sec_clk_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17512\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22225\,
            ce => 'H',
            sr => \N__20681\
        );

    \CONSTANT_ONE_LUT4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => \CONSTANT_ONE_NET_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001101011010"
        )
    port map (
            in0 => \N__9726\,
            in1 => \N__9859\,
            in2 => \N__9291\,
            in3 => \N__9536\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22217\,
            ce => \N__9652\,
            sr => \N__20683\
        );

    \buart.Z_rx.bitcount_es_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__9858\,
            in1 => \N__9288\,
            in2 => \N__9545\,
            in3 => \N__9279\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22217\,
            ce => \N__9652\,
            sr => \N__20683\
        );

    \uu0.delay_line_RNILLLG7_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__9249\,
            in1 => \N__9240\,
            in2 => \_gnd_net_\,
            in3 => \N__9225\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16245\,
            in1 => \N__12111\,
            in2 => \_gnd_net_\,
            in3 => \N__21772\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13016\,
            in1 => \N__9567\,
            in2 => \_gnd_net_\,
            in3 => \N__9667\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14961\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9489\,
            lcout => \resetGen.un241_ci\,
            ltout => \resetGen.un241_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011010"
        )
    port map (
            in0 => \N__9462\,
            in1 => \N__9438\,
            in2 => \N__9513\,
            in3 => \N__11175\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9509\,
            in1 => \N__9490\,
            in2 => \_gnd_net_\,
            in3 => \N__9461\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011010"
        )
    port map (
            in0 => \N__9471\,
            in1 => \N__9439\,
            in2 => \N__9474\,
            in3 => \N__11176\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9470\,
            in2 => \_gnd_net_\,
            in3 => \N__9460\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__9450\,
            in1 => \N__9437\,
            in2 => \N__9444\,
            in3 => \N__11177\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9735\,
            in1 => \N__9882\,
            in2 => \_gnd_net_\,
            in3 => \N__9725\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9847\,
            in2 => \_gnd_net_\,
            in3 => \N__9598\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9910\,
            in1 => \N__9933\,
            in2 => \N__9800\,
            in3 => \N__9619\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9958\,
            in2 => \N__9678\,
            in3 => \N__9597\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__9846\,
            in1 => \N__9942\,
            in2 => \N__9675\,
            in3 => \N__9960\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__9884\,
            in1 => \N__9848\,
            in2 => \N__9915\,
            in3 => \N__9894\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9845\,
            in1 => \_gnd_net_\,
            in2 => \N__9605\,
            in3 => \N__9620\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__9883\,
            in1 => \N__9844\,
            in2 => \N__9672\,
            in3 => \N__14962\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9621\,
            in2 => \N__9606\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9959\,
            in2 => \_gnd_net_\,
            in3 => \N__9936\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9866\,
            in1 => \N__9932\,
            in2 => \_gnd_net_\,
            in3 => \N__9918\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__22197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9911\,
            in2 => \_gnd_net_\,
            in3 => \N__9888\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__9885\,
            in1 => \N__9865\,
            in2 => \N__9801\,
            in3 => \N__9804\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_3_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10274\,
            in1 => \N__10243\,
            in2 => \N__9758\,
            in3 => \N__10214\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__10182\,
            sr => \N__20674\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10477\,
            in2 => \_gnd_net_\,
            in3 => \N__10113\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9776\,
            in1 => \N__10005\,
            in2 => \N__9783\,
            in3 => \N__10068\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__10182\,
            sr => \N__20674\
        );

    \uu2.r_addr_esr_7_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10069\,
            in1 => \N__10046\,
            in2 => \N__10028\,
            in3 => \N__9765\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__10182\,
            sr => \N__20674\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10273\,
            in1 => \N__10242\,
            in2 => \N__9757\,
            in3 => \N__10213\,
            lcout => \uu2.un404_ci_0\,
            ltout => \uu2.un404_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__10024\,
            in1 => \N__10478\,
            in2 => \N__10053\,
            in3 => \N__10114\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__10182\,
            sr => \N__20674\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10045\,
            in2 => \_gnd_net_\,
            in3 => \N__10020\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__13197\,
            in1 => \N__13304\,
            in2 => \N__13431\,
            in3 => \N__13384\,
            lcout => \uu2.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__21766\,
            in1 => \N__12993\,
            in2 => \N__11319\,
            in3 => \N__11127\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__9987\,
            in1 => \N__10965\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__11291\,
            in1 => \N__11311\,
            in2 => \_gnd_net_\,
            in3 => \N__12991\,
            lcout => \uu2.N_34\,
            ltout => \uu2.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__10905\,
            in1 => \N__21768\,
            in2 => \N__9981\,
            in3 => \N__10700\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__10701\,
            in1 => \N__10293\,
            in2 => \N__21787\,
            in3 => \N__11022\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__10842\,
            in2 => \_gnd_net_\,
            in3 => \N__21764\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__11292\,
            in1 => \N__12992\,
            in2 => \N__11318\,
            in3 => \N__12107\,
            lcout => \uu2.N_31\,
            ltout => \uu2.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21767\,
            in2 => \N__10284\,
            in3 => \N__10884\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_2_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10142\,
            in1 => \N__10269\,
            in2 => \N__10247\,
            in3 => \N__10209\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22253\,
            ce => 'H',
            sr => \N__20668\
        );

    \uu2.r_addr_1_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10208\,
            in1 => \N__10238\,
            in2 => \_gnd_net_\,
            in3 => \N__10140\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22253\,
            ce => 'H',
            sr => \N__20668\
        );

    \uu2.r_addr_0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10207\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22253\,
            ce => 'H',
            sr => \N__20668\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10138\,
            in2 => \_gnd_net_\,
            in3 => \N__20761\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_4_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10106\,
            in1 => \N__10076\,
            in2 => \_gnd_net_\,
            in3 => \N__10141\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22253\,
            ce => 'H',
            sr => \N__20668\
        );

    \uu2.vram_rd_clk_det_0_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10170\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.vram_rd_clk_det_0C_net\,
            ce => 'H',
            sr => \N__20629\
        );

    \uu2.r_addr_5_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10146\,
            in1 => \N__10115\,
            in2 => \N__10476\,
            in3 => \N__10080\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22238\,
            ce => 'H',
            sr => \N__20661\
        );

    \uu2.l_count_7_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10446\,
            in1 => \N__10363\,
            in2 => \N__10419\,
            in3 => \N__10398\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22238\,
            ce => 'H',
            sr => \N__20661\
        );

    \Lab_UT.didp.reset_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11436\,
            in1 => \_gnd_net_\,
            in2 => \N__12279\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22238\,
            ce => 'H',
            sr => \N__20661\
        );

    \Lab_UT.didp.ce_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12275\,
            in2 => \_gnd_net_\,
            in3 => \N__11435\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22238\,
            ce => 'H',
            sr => \N__20661\
        );

    \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14811\,
            in2 => \_gnd_net_\,
            in3 => \N__20754\,
            lcout => \Lab_UT.didp.regrce3.LdAMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10311\,
            in2 => \_gnd_net_\,
            in3 => \N__10617\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__10618\,
            in1 => \_gnd_net_\,
            in2 => \N__10323\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22238\,
            ce => 'H',
            sr => \N__20661\
        );

    \Lab_UT.didp.regrce4.q_esr_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20050\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => \N__10986\,
            sr => \N__20659\
        );

    \Lab_UT.didp.regrce4.q_esr_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21390\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => \N__10986\,
            sr => \N__20659\
        );

    \Lab_UT.didp.regrce4.q_esr_2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20956\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => \N__10986\,
            sr => \N__20659\
        );

    \Lab_UT.didp.regrce4.q_esr_3_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21140\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => \N__10986\,
            sr => \N__20659\
        );

    \uu2.vram_wr_en_0_i_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111110101111"
        )
    port map (
            in0 => \N__10796\,
            in1 => \N__10943\,
            in2 => \N__22281\,
            in3 => \N__10863\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__14293\,
            in1 => \N__20046\,
            in2 => \_gnd_net_\,
            in3 => \N__14361\,
            lcout => \Lab_UT.didp.countrce1.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_3_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__11048\,
            in1 => \N__10497\,
            in2 => \N__11096\,
            in3 => \N__10488\,
            lcout => \G_188\,
            ltout => \G_188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__18119\,
            in1 => \N__11587\,
            in2 => \N__10491\,
            in3 => \N__11460\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101000101"
        )
    port map (
            in0 => \N__10821\,
            in1 => \N__10658\,
            in2 => \N__11592\,
            in3 => \N__18121\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_armed_2_0_iso_i_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11693\,
            in2 => \_gnd_net_\,
            in3 => \N__11646\,
            lcout => \Lab_UT.un1_armed_2_0_iso_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_rst_0_iclk_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__20749\,
            in1 => \_gnd_net_\,
            in2 => \N__11708\,
            in3 => \N__11647\,
            lcout => \Lab_UT.un1_rst_0_iclkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__10820\,
            in1 => \N__10657\,
            in2 => \N__11591\,
            in3 => \N__18120\,
            lcout => \Lab_UT.dispString.dOutP_1_iv_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11701\,
            in2 => \_gnd_net_\,
            in3 => \N__11650\,
            lcout => \G_182\,
            ltout => \G_182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_4_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__11702\,
            in1 => \N__20755\,
            in2 => \N__10662\,
            in3 => \N__10659\,
            lcout => \G_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__10641\,
            in1 => \N__11495\,
            in2 => \N__11769\,
            in3 => \N__10629\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.justentered_latch_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__11494\,
            in1 => \N__10639\,
            in2 => \N__10644\,
            in3 => \N__20756\,
            lcout => \G_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__10640\,
            in1 => \N__10628\,
            in2 => \N__11768\,
            in3 => \N__11493\,
            lcout => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10599\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22198\,
            ce => 'H',
            sr => \N__20688\
        );

    \buart.Z_tx.shifter_7_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20451\,
            in1 => \N__10539\,
            in2 => \_gnd_net_\,
            in3 => \N__10572\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22259\,
            ce => \N__20372\,
            sr => \N__20693\
        );

    \buart.Z_tx.shifter_8_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20452\,
            in2 => \_gnd_net_\,
            in3 => \N__10548\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22259\,
            ce => \N__20372\,
            sr => \N__20693\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15978\,
            in1 => \N__21748\,
            in2 => \_gnd_net_\,
            in3 => \N__13262\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10734\,
            in1 => \N__10719\,
            in2 => \_gnd_net_\,
            in3 => \N__20747\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__21692\,
            in1 => \N__20273\,
            in2 => \_gnd_net_\,
            in3 => \N__13383\,
            lcout => \uu2.w_addr_displaying_RNI03P31Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__16260\,
            in1 => \N__10797\,
            in2 => \_gnd_net_\,
            in3 => \N__10809\,
            lcout => \uu2.un28_w_addr_user_i\,
            ltout => \uu2.un28_w_addr_user_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNID65PE_4_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10671\,
            in3 => \N__15929\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI43E87_4_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__16259\,
            in1 => \N__20746\,
            in2 => \_gnd_net_\,
            in3 => \N__10808\,
            lcout => \uu2.w_addr_user_RNI43E87Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000111011110"
        )
    port map (
            in0 => \N__16554\,
            in1 => \N__13386\,
            in2 => \N__13789\,
            in3 => \N__12137\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101000010"
        )
    port map (
            in0 => \N__12106\,
            in1 => \N__16106\,
            in2 => \N__10668\,
            in3 => \N__11279\,
            lcout => \uu2.bitmap_pmux_sn_i5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11388\,
            in2 => \_gnd_net_\,
            in3 => \N__13385\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010010"
        )
    port map (
            in0 => \N__12138\,
            in1 => \N__16623\,
            in2 => \N__11397\,
            in3 => \N__13782\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13743\,
            in2 => \N__10665\,
            in3 => \N__11952\,
            lcout => \uu2.N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16555\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__11901\,
            sr => \N__20617\
        );

    \uu2.w_addr_displaying_fast_nesr_1_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11393\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__11901\,
            sr => \N__20617\
        );

    \uu2.w_addr_displaying_nesr_1_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16557\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__11901\,
            sr => \N__20617\
        );

    \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10686\,
            in1 => \N__10740\,
            in2 => \_gnd_net_\,
            in3 => \N__10710\,
            lcout => OPEN,
            ltout => \uu2.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__11256\,
            in1 => \N__10764\,
            in2 => \N__10704\,
            in3 => \N__11325\,
            lcout => \uu2.bitmap_pmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__13777\,
            in1 => \N__13263\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNICM7R_180_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16371\,
            in1 => \N__12243\,
            in2 => \_gnd_net_\,
            in3 => \N__11936\,
            lcout => OPEN,
            ltout => \uu2.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__13778\,
            in1 => \N__16631\,
            in2 => \N__10692\,
            in3 => \N__12219\,
            lcout => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\,
            ltout => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__12005\,
            in1 => \N__10757\,
            in2 => \N__10689\,
            in3 => \N__16313\,
            lcout => \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__13264\,
            in1 => \N__10770\,
            in2 => \_gnd_net_\,
            in3 => \N__16632\,
            lcout => \uu2.bitmap_pmux_u_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__10758\,
            in1 => \N__16314\,
            in2 => \N__12009\,
            in3 => \N__10746\,
            lcout => \uu2.w_addr_displaying_RNI0NG56Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_1_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10733\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.vram_rd_clk_det_1C_net\,
            ce => 'H',
            sr => \N__20630\
        );

    \Lab_UT.didp.regrce3.q_esr_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20052\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22232\,
            ce => \N__14621\,
            sr => \N__20664\
        );

    \Lab_UT.didp.regrce3.q_esr_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20945\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22232\,
            ce => \N__14621\,
            sr => \N__20664\
        );

    \Lab_UT.didp.regrce3.q_esr_3_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21121\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22232\,
            ce => \N__14621\,
            sr => \N__20664\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__18002\,
            in1 => \N__17123\,
            in2 => \N__11523\,
            in3 => \N__13612\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_1_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18201\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22226\,
            ce => 'H',
            sr => \N__20662\
        );

    \Lab_UT.dispString.cnt_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__18003\,
            in1 => \N__17492\,
            in2 => \N__18220\,
            in3 => \N__18081\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22226\,
            ce => 'H',
            sr => \N__20662\
        );

    \Lab_UT.didp.ce_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17491\,
            in1 => \N__12687\,
            in2 => \_gnd_net_\,
            in3 => \N__18478\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22226\,
            ce => 'H',
            sr => \N__20662\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__14420\,
            in1 => \N__12173\,
            in2 => \N__14546\,
            in3 => \N__17122\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12564\,
            in2 => \N__10812\,
            in3 => \N__14680\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17294\,
            in1 => \N__13579\,
            in2 => \N__17087\,
            in3 => \N__12517\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_0_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__10862\,
            in1 => \_gnd_net_\,
            in2 => \N__10944\,
            in3 => \N__10792\,
            lcout => \uu2.un4_w_user_data_rdyZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un20_w_addr_user_1_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__10911\,
            in1 => \N__10939\,
            in2 => \N__10974\,
            in3 => \N__10861\,
            lcout => \uu2.un20_w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18197\,
            in1 => \N__18007\,
            in2 => \N__17493\,
            in3 => \N__18079\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18078\,
            in1 => \N__18196\,
            in2 => \_gnd_net_\,
            in3 => \N__11148\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__14547\,
            in1 => \N__12495\,
            in2 => \N__10776\,
            in3 => \N__12401\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__17429\,
            in1 => \N__11552\,
            in2 => \N__10773\,
            in3 => \N__13650\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__19137\,
            in1 => \N__18477\,
            in2 => \N__20766\,
            in3 => \N__19511\,
            lcout => \Lab_UT.didp.regrce4.LdAMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__10835\,
            in2 => \N__10964\,
            in3 => \N__11012\,
            lcout => \uu2.un1_w_user_lfZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__18115\,
            in1 => \N__11146\,
            in2 => \N__17430\,
            in3 => \N__11581\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_4_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10957\,
            in1 => \N__21869\,
            in2 => \N__11123\,
            in3 => \N__11011\,
            lcout => \uu2.un1_w_user_crZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__11551\,
            in1 => \N__10926\,
            in2 => \N__13686\,
            in3 => \N__10917\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_3_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10898\,
            in1 => \N__11116\,
            in2 => \_gnd_net_\,
            in3 => \N__21868\,
            lcout => \uu2.un1_w_user_lfZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_3_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10834\,
            in1 => \N__10897\,
            in2 => \_gnd_net_\,
            in3 => \N__10876\,
            lcout => \uu2.un1_w_user_crZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__18012\,
            in1 => \N__18116\,
            in2 => \_gnd_net_\,
            in3 => \N__10848\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIKUO21_1_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__18226\,
            in1 => \N__17542\,
            in2 => \N__17571\,
            in3 => \N__12542\,
            lcout => \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101010101"
        )
    port map (
            in0 => \N__11651\,
            in1 => \N__11147\,
            in2 => \N__20765\,
            in3 => \N__11703\,
            lcout => \G_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18123\,
            in1 => \N__11583\,
            in2 => \_gnd_net_\,
            in3 => \N__11198\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_idle_4_0_iclk_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__11704\,
            in1 => \N__11652\,
            in2 => \_gnd_net_\,
            in3 => \N__11215\,
            lcout => OPEN,
            ltout => \Lab_UT.un1_idle_4_0_iclkZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_1_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__11094\,
            in1 => \N__11049\,
            in2 => \N__11037\,
            in3 => \N__11034\,
            lcout => \G_185\,
            ltout => \G_185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11582\,
            in2 => \N__11028\,
            in3 => \N__18122\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__11544\,
            in1 => \N__11409\,
            in2 => \N__11025\,
            in3 => \N__17831\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__20764\,
            in1 => \N__11699\,
            in2 => \_gnd_net_\,
            in3 => \N__11654\,
            lcout => \G_180\,
            ltout => \G_180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__11700\,
            in1 => \N__10998\,
            in2 => \N__10992\,
            in3 => \N__11217\,
            lcout => \G_181\,
            ltout => \G_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_0__m3_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__11496\,
            in1 => \N__11653\,
            in2 => \N__10989\,
            in3 => \N__11753\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__11655\,
            in1 => \N__11226\,
            in2 => \N__11220\,
            in3 => \N__11216\,
            lcout => \G_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m59_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11648\,
            in1 => \N__14910\,
            in2 => \_gnd_net_\,
            in3 => \N__11697\,
            lcout => \Lab_UT.alarmstate_0_sqmuxa_1\,
            ltout => \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_6_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000110"
        )
    port map (
            in0 => \N__11698\,
            in1 => \N__11649\,
            in2 => \N__11202\,
            in3 => \N__11199\,
            lcout => \G_184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m37_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12906\,
            in1 => \N__13091\,
            in2 => \N__11742\,
            in3 => \N__12811\,
            lcout => \Lab_UT.dictrl.next_state6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13093\,
            in1 => \N__15747\,
            in2 => \N__20928\,
            in3 => \N__12812\,
            lcout => OPEN,
            ltout => \resetGen.escKeyZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11154\,
            in2 => \N__11187\,
            in3 => \N__14974\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_4_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21313\,
            in1 => \N__19990\,
            in2 => \N__15610\,
            in3 => \N__21097\,
            lcout => \resetGen.escKeyZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__21312\,
            in2 => \_gnd_net_\,
            in3 => \N__20904\,
            lcout => \Lab_UT.dictrl.g2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_5_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__13092\,
            in1 => \N__15746\,
            in2 => \N__18479\,
            in3 => \N__15596\,
            lcout => \Lab_UT.dictrl.G_25_i_o3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21306\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22193\,
            ce => \N__20794\,
            sr => \N__20690\
        );

    \buart.Z_rx.shifter_1_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20900\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22193\,
            ce => \N__20794\,
            sr => \N__20690\
        );

    \buart.Z_rx.shifter_3_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15602\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22193\,
            ce => \N__20794\,
            sr => \N__20690\
        );

    \buart.Z_rx.shifter_7_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13028\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22190\,
            ce => \N__20792\,
            sr => \N__20692\
        );

    \uu2.w_addr_user_2_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__21836\,
            in1 => \N__16231\,
            in2 => \N__20341\,
            in3 => \N__11245\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_user_1_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__11243\,
            in1 => \_gnd_net_\,
            in2 => \N__16238\,
            in3 => \N__20332\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_user_0_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16227\,
            in2 => \_gnd_net_\,
            in3 => \N__11242\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_user_4_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11244\,
            in1 => \N__16012\,
            in2 => \_gnd_net_\,
            in3 => \N__16294\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_user_5_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16295\,
            in1 => \N__15521\,
            in2 => \N__16017\,
            in3 => \N__11246\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_user_6_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11247\,
            in1 => \N__16016\,
            in2 => \N__16039\,
            in3 => \N__16193\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15941\
        );

    \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20748\,
            in2 => \_gnd_net_\,
            in3 => \N__15879\,
            lcout => \uu2.N_33_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIKIPH1_8_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20275\,
            in1 => \N__21676\,
            in2 => \N__16121\,
            in3 => \N__13266\,
            lcout => \uu2.un51_w_data_displaying_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12079\,
            in2 => \_gnd_net_\,
            in3 => \N__20274\,
            lcout => OPEN,
            ltout => \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIASLS1_8_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21675\,
            in1 => \N__16113\,
            in2 => \N__11295\,
            in3 => \N__13265\,
            lcout => \uu2.w_data_displaying_2_i_a2_i_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_3_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16114\,
            in1 => \N__20278\,
            in2 => \N__21688\,
            in3 => \N__12084\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__11890\,
            sr => \N__20620\
        );

    \uu2.w_addr_displaying_fast_nesr_3_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20276\,
            in1 => \N__21678\,
            in2 => \N__12099\,
            in3 => \N__11937\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__11890\,
            sr => \N__20620\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21677\,
            in1 => \N__20277\,
            in2 => \N__13790\,
            in3 => \N__12080\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__11890\,
            sr => \N__20620\
        );

    \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001000"
        )
    port map (
            in0 => \N__21674\,
            in1 => \N__13161\,
            in2 => \N__16120\,
            in3 => \N__11280\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0FGN6_4_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11268\,
            in2 => \N__11259\,
            in3 => \N__12015\,
            lcout => \uu2.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__16482\,
            in1 => \N__16451\,
            in2 => \N__17724\,
            in3 => \N__16920\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__20618\
        );

    \uu2.bitmap_221_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__16919\,
            in1 => \N__17720\,
            in2 => \N__16452\,
            in3 => \N__16481\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__20618\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16542\,
            in2 => \_gnd_net_\,
            in3 => \N__11396\,
            lcout => \uu2.N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIPIHG1_75_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__16543\,
            in1 => \N__11991\,
            in2 => \N__11985\,
            in3 => \N__14001\,
            lcout => OPEN,
            ltout => \uu2.N_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__16116\,
            in1 => \N__11345\,
            in2 => \N__11364\,
            in3 => \N__12192\,
            lcout => \uu2.bitmap_pmux_27_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI6MCU1_93_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__16544\,
            in1 => \N__11361\,
            in2 => \N__11355\,
            in3 => \N__16491\,
            lcout => OPEN,
            ltout => \uu2.N_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI72CH8_69_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__11346\,
            in1 => \N__11907\,
            in2 => \N__11334\,
            in3 => \N__11331\,
            lcout => \uu2.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_3_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12273\,
            in1 => \N__14186\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__20669\
        );

    \Lab_UT.didp.ce_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12185\,
            in1 => \N__17884\,
            in2 => \N__17496\,
            in3 => \N__13726\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__20669\
        );

    \Lab_UT.didp.reset_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__13727\,
            in1 => \N__17487\,
            in2 => \N__17891\,
            in3 => \N__12186\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__20669\
        );

    \Lab_UT.didp.reset_2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12274\,
            in1 => \N__14187\,
            in2 => \_gnd_net_\,
            in3 => \N__11429\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__20669\
        );

    \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12184\,
            in1 => \N__17883\,
            in2 => \N__17495\,
            in3 => \N__13725\,
            lcout => \Lab_UT.didp.ce_12_1\,
            ltout => \Lab_UT.didp.ce_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12262\,
            in2 => \N__11415\,
            in3 => \N__14185\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16758\,
            in1 => \N__17619\,
            in2 => \N__11412\,
            in3 => \N__13508\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__20669\
        );

    \Lab_UT.didp.countrce2.q_3_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__12482\,
            in1 => \N__12327\,
            in2 => \N__12465\,
            in3 => \N__12305\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001011"
        )
    port map (
            in0 => \N__13854\,
            in1 => \N__12483\,
            in2 => \N__12321\,
            in3 => \N__12459\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__16749\,
            in1 => \N__12397\,
            in2 => \N__12626\,
            in3 => \N__12169\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13853\,
            in1 => \N__12364\,
            in2 => \N__12309\,
            in3 => \N__14579\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__14559\,
            in1 => \N__12559\,
            in2 => \N__17494\,
            in3 => \N__14519\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17877\,
            in1 => \N__14346\,
            in2 => \_gnd_net_\,
            in3 => \N__16989\,
            lcout => \Lab_UT.didp.countrce1.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__18194\,
            in1 => \N__18077\,
            in2 => \N__18008\,
            in3 => \N__12365\,
            lcout => \Lab_UT.dispString.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13491\,
            in1 => \N__13675\,
            in2 => \N__13721\,
            in3 => \N__13534\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12336\,
            in1 => \N__14172\,
            in2 => \N__11514\,
            in3 => \N__11511\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11505\,
            in1 => \N__12408\,
            in2 => \N__11499\,
            in3 => \N__11442\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__13709\,
            in1 => \N__14292\,
            in2 => \N__11472\,
            in3 => \N__21116\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__14251\,
            in1 => \N__14210\,
            in2 => \N__11463\,
            in3 => \N__13710\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_3_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__18195\,
            in1 => \N__12558\,
            in2 => \N__17480\,
            in3 => \N__13535\,
            lcout => \Lab_UT.dispString.N_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__13631\,
            in1 => \N__14336\,
            in2 => \N__11601\,
            in3 => \N__11448\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17679\,
            in1 => \N__21117\,
            in2 => \N__12153\,
            in3 => \N__13497\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__13498\,
            in1 => \N__16831\,
            in2 => \N__11730\,
            in3 => \N__16788\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__11727\,
            in1 => \N__16942\,
            in2 => \N__11553\,
            in3 => \N__11718\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__17677\,
            in1 => \N__20031\,
            in2 => \_gnd_net_\,
            in3 => \N__17083\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000001"
        )
    port map (
            in0 => \N__16830\,
            in1 => \N__16808\,
            in2 => \N__11712\,
            in3 => \N__17678\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__13619\,
            in1 => \N__16707\,
            in2 => \N__11709\,
            in3 => \N__11645\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIH15E_2_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17982\,
            in2 => \_gnd_net_\,
            in3 => \N__18228\,
            lcout => \Lab_UT.dispString.un42_dOutP_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIOG7L_2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__18114\,
            in1 => \N__17997\,
            in2 => \_gnd_net_\,
            in3 => \N__18227\,
            lcout => \Lab_UT.dispString.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17981\,
            in2 => \_gnd_net_\,
            in3 => \N__18113\,
            lcout => \Lab_UT.dispString.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14844\,
            in2 => \_gnd_net_\,
            in3 => \N__20762\,
            lcout => \Lab_UT.didp.regrce2.LdAStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20032\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22196\,
            ce => \N__11778\,
            sr => \N__20665\
        );

    \Lab_UT.didp.regrce2.q_esr_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21352\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22196\,
            ce => \N__11778\,
            sr => \N__20665\
        );

    \Lab_UT.didp.regrce2.q_esr_2_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22196\,
            ce => \N__11778\,
            sr => \N__20665\
        );

    \Lab_UT.didp.regrce2.q_esr_3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21094\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22196\,
            ce => \N__11778\,
            sr => \N__20665\
        );

    \Lab_UT.dictrl.alarmstate8_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13103\,
            in1 => \N__15741\,
            in2 => \N__19036\,
            in3 => \N__11784\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_5_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15743\,
            in1 => \N__12823\,
            in2 => \N__19774\,
            in3 => \N__15609\,
            lcout => \Lab_UT.dictrl.g1_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m37_N_2L1_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20006\,
            in1 => \N__15742\,
            in2 => \N__20927\,
            in3 => \N__21231\,
            lcout => \Lab_UT.dictrl.m37_N_2LZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__12824\,
            in1 => \N__21092\,
            in2 => \N__13112\,
            in3 => \N__15744\,
            lcout => \Lab_UT.dictrl.g0_5_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21232\,
            in1 => \N__13104\,
            in2 => \_gnd_net_\,
            in3 => \N__19696\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__17239\,
            in1 => \N__11814\,
            in2 => \N__11808\,
            in3 => \N__21336\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__11805\,
            in1 => \N__11793\,
            in2 => \N__11799\,
            in3 => \N__19923\,
            lcout => \Lab_UT.dictrl.N_55_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_6_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15745\,
            in2 => \_gnd_net_\,
            in3 => \N__12807\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19510\,
            in1 => \N__15587\,
            in2 => \N__11796\,
            in3 => \N__13101\,
            lcout => \Lab_UT.dictrl.g0_6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__20908\,
            in1 => \N__19509\,
            in2 => \N__15603\,
            in3 => \N__21314\,
            lcout => \Lab_UT.dictrl.g0_5_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111111"
        )
    port map (
            in0 => \N__12808\,
            in1 => \_gnd_net_\,
            in2 => \N__19929\,
            in3 => \N__20139\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_25_i_o3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__21054\,
            in1 => \N__21315\,
            in2 => \N__11787\,
            in3 => \N__20909\,
            lcout => \Lab_UT.dictrl.G_25_i_o3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_3_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15583\,
            in1 => \N__12806\,
            in2 => \N__21213\,
            in3 => \N__19668\,
            lcout => \Lab_UT.dictrl.alarmstate8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21307\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_6_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13102\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_fast_4_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15739\,
            lcout => \buart__rx_shifter_fast_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_0_rep1_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21308\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_fast_2_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21044\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_3_rep2_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15600\,
            lcout => bu_rx_data_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15738\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => \N__20795\,
            sr => \N__20691\
        );

    \buart.Z_rx.shifter_2_rep1_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21084\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22189\,
            ce => \N__20793\,
            sr => \N__20694\
        );

    \buart.Z_rx.shifter_5_rep1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22189\,
            ce => \N__20793\,
            sr => \N__20694\
        );

    \buart.Z_rx.shifter_fast_5_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12821\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22189\,
            ce => \N__20793\,
            sr => \N__20694\
        );

    \buart.Z_rx.shifter_fast_3_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15601\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22189\,
            ce => \N__20793\,
            sr => \N__20694\
        );

    \buart.Z_rx.shifter_5_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12825\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22188\,
            ce => \N__20790\,
            sr => \N__20695\
        );

    \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__16633\,
            in1 => \N__13296\,
            in2 => \N__13193\,
            in3 => \N__13369\,
            lcout => \uu2.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_6_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101111000011"
        )
    port map (
            in0 => \N__13249\,
            in1 => \N__13189\,
            in2 => \N__13323\,
            in3 => \N__16635\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_ness_6C_net\,
            ce => \N__11897\,
            sr => \N__20624\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__13188\,
            in1 => \_gnd_net_\,
            in2 => \N__21803\,
            in3 => \N__16181\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13370\,
            in1 => \N__16289\,
            in2 => \_gnd_net_\,
            in3 => \N__21788\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21789\,
            in1 => \N__15519\,
            in2 => \_gnd_net_\,
            in3 => \N__13297\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16290\,
            lcout => \uu2.un426_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__16634\,
            in1 => \_gnd_net_\,
            in2 => \N__21804\,
            in3 => \N__16160\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16191\,
            lcout => \uu2.vbuf_w_addr_user.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_168_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__13908\,
            in1 => \N__14151\,
            in2 => \N__13946\,
            in3 => \N__13974\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__20623\
        );

    \uu2.bitmap_40_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__13976\,
            in1 => \N__13941\,
            in2 => \N__14160\,
            in3 => \N__13910\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__20623\
        );

    \uu2.bitmap_75_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__13911\,
            in1 => \N__14158\,
            in2 => \N__13947\,
            in3 => \N__13977\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__20623\
        );

    \uu2.bitmap_203_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__13975\,
            in1 => \N__13940\,
            in2 => \N__14159\,
            in3 => \N__13909\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__20623\
        );

    \uu2.bitmap_RNIJS4P_162_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11933\,
            in1 => \N__11976\,
            in2 => \_gnd_net_\,
            in3 => \N__13131\,
            lcout => \uu2.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__12127\,
            in1 => \N__11970\,
            in2 => \_gnd_net_\,
            in3 => \N__11935\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16647\,
            in2 => \N__11961\,
            in3 => \N__11958\,
            lcout => \uu2.bitmap_RNI2Q8F1Z0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIBPBO_40_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111000111"
        )
    port map (
            in0 => \N__11943\,
            in1 => \N__11934\,
            in2 => \N__16353\,
            in3 => \N__13881\,
            lcout => \uu2.bitmap_pmux_26_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_197_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__13563\,
            in1 => \N__14664\,
            in2 => \N__13473\,
            in3 => \N__14490\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20621\
        );

    \uu2.bitmap_RNITSCU1_69_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__13137\,
            in1 => \N__11913\,
            in2 => \N__12093\,
            in3 => \N__13734\,
            lcout => \uu2.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12072\,
            in2 => \_gnd_net_\,
            in3 => \N__15889\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20621\
        );

    \uu2.w_addr_displaying_fast_2_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15891\,
            in1 => \N__20297\,
            in2 => \N__12095\,
            in3 => \N__12131\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20621\
        );

    \uu2.w_addr_displaying_2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__15890\,
            in2 => \N__12092\,
            in3 => \N__21673\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20621\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21672\,
            in1 => \N__16099\,
            in2 => \N__12094\,
            in3 => \N__20295\,
            lcout => \uu2.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000100000000"
        )
    port map (
            in0 => \N__16098\,
            in1 => \N__21671\,
            in2 => \N__12091\,
            in3 => \N__13314\,
            lcout => \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIGEPH1_4_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101000001000"
        )
    port map (
            in0 => \N__21670\,
            in1 => \N__20294\,
            in2 => \N__16115\,
            in3 => \N__13382\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100011001"
        )
    port map (
            in0 => \N__14060\,
            in1 => \N__14388\,
            in2 => \N__14111\,
            in3 => \N__13830\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_212_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__14387\,
            in1 => \N__13829\,
            in2 => \N__14110\,
            in3 => \N__14059\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_84_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000111101"
        )
    port map (
            in0 => \N__14062\,
            in1 => \N__14390\,
            in2 => \N__14113\,
            in3 => \N__13832\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_180_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__14386\,
            in1 => \N__13828\,
            in2 => \N__14109\,
            in3 => \N__14058\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_52_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111101111001"
        )
    port map (
            in0 => \N__14061\,
            in1 => \N__14389\,
            in2 => \N__14112\,
            in3 => \N__13831\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_RNIB3QK_52_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16349\,
            in1 => \N__12231\,
            in2 => \_gnd_net_\,
            in3 => \N__12225\,
            lcout => \uu2.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__14063\,
            in1 => \N__14391\,
            in2 => \N__14114\,
            in3 => \N__13833\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20619\
        );

    \uu2.bitmap_RNIRMQA1_84_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__12207\,
            in1 => \N__16407\,
            in2 => \N__12201\,
            in3 => \N__14025\,
            lcout => \uu2.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17790\,
            in1 => \N__17301\,
            in2 => \_gnd_net_\,
            in3 => \N__12518\,
            lcout => \Lab_UT.min2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14355\,
            in2 => \_gnd_net_\,
            in3 => \N__16979\,
            lcout => \Lab_UT.didp.countrce1.ce_12_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17791\,
            in1 => \N__16747\,
            in2 => \_gnd_net_\,
            in3 => \N__12174\,
            lcout => \Lab_UT.min2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17037\,
            in1 => \N__17618\,
            in2 => \_gnd_net_\,
            in3 => \N__17101\,
            lcout => \Lab_UT.didp.countrce4.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_2_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12627\,
            in3 => \N__13865\,
            lcout => \Lab_UT.didp.countrce2.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17792\,
            in1 => \N__12620\,
            in2 => \_gnd_net_\,
            in3 => \N__12402\,
            lcout => \Lab_UT.sec1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12372\,
            in1 => \N__12306\,
            in2 => \_gnd_net_\,
            in3 => \N__17793\,
            lcout => \Lab_UT.sec1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__14454\,
            in1 => \N__12655\,
            in2 => \N__12345\,
            in3 => \N__20946\,
            lcout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17029\,
            in1 => \N__16943\,
            in2 => \N__16985\,
            in3 => \N__14515\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__14453\,
            in1 => \_gnd_net_\,
            in2 => \N__12625\,
            in3 => \N__13870\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__12656\,
            in1 => \N__12308\,
            in2 => \N__12330\,
            in3 => \N__21136\,
            lcout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100001111"
        )
    port map (
            in0 => \N__12615\,
            in1 => \N__13871\,
            in2 => \N__21391\,
            in3 => \N__12657\,
            lcout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18473\,
            in1 => \N__19922\,
            in2 => \N__17252\,
            in3 => \N__18346\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14452\,
            in1 => \N__12307\,
            in2 => \N__12624\,
            in3 => \N__13869\,
            lcout => \Lab_UT.didp.un24_ce_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__17124\,
            in1 => \N__13589\,
            in2 => \N__12563\,
            in3 => \N__12522\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI62AM_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12431\,
            in2 => \_gnd_net_\,
            in3 => \N__12646\,
            lcout => \Lab_UT.didp.un1_dicLdStens_0\,
            ltout => \Lab_UT.didp.un1_dicLdStens_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__14439\,
            in1 => \N__12474\,
            in2 => \N__12468\,
            in3 => \N__12464\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101000001"
        )
    port map (
            in0 => \N__12463\,
            in1 => \N__12647\,
            in2 => \N__12579\,
            in3 => \N__12432\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__14208\,
            in1 => \N__12420\,
            in2 => \N__14258\,
            in3 => \N__14351\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17036\,
            in2 => \_gnd_net_\,
            in3 => \N__17077\,
            lcout => \Lab_UT.didp.countrce4.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__14410\,
            in2 => \N__14450\,
            in3 => \N__17827\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20757\,
            in2 => \_gnd_net_\,
            in3 => \N__18246\,
            lcout => \Lab_UT.didp.regrce1.LdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__17866\,
            in1 => \N__14209\,
            in2 => \N__14259\,
            in3 => \N__12570\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_esr_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15069\,
            in1 => \N__18603\,
            in2 => \N__15224\,
            in3 => \N__15029\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => \N__18514\,
            sr => \N__20660\
        );

    \Lab_UT.dictrl.state_ret_11_ess_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__15030\,
            in1 => \N__15220\,
            in2 => \N__18611\,
            in3 => \N__15070\,
            lcout => \Lab_UT.LdSones_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => \N__18514\,
            sr => \N__20660\
        );

    \Lab_UT.dictrl.state_ret_8_ess_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__15071\,
            in1 => \N__18607\,
            in2 => \N__15225\,
            in3 => \N__15031\,
            lcout => \Lab_UT.state_ret_8_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => \N__18514\,
            sr => \N__20660\
        );

    \Lab_UT.didp.state_ret_1_esr_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__15032\,
            in1 => \_gnd_net_\,
            in2 => \N__18612\,
            in3 => \N__15072\,
            lcout => \Lab_UT.didp.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => \N__18514\,
            sr => \N__20660\
        );

    \Lab_UT.didp.ce_RNIFQ9K_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12675\,
            in2 => \_gnd_net_\,
            in3 => \N__12669\,
            lcout => \Lab_UT.didp.un1_dicLdSones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__12645\,
            in1 => \N__20030\,
            in2 => \_gnd_net_\,
            in3 => \N__12616\,
            lcout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__21377\,
            in1 => \N__14347\,
            in2 => \N__14294\,
            in3 => \N__17881\,
            lcout => \Lab_UT.didp.countrce1.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22205\,
            ce => \N__12705\,
            sr => \N__20666\
        );

    \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20958\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22205\,
            ce => \N__12705\,
            sr => \N__20666\
        );

    \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21141\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22205\,
            ce => \N__12705\,
            sr => \N__20666\
        );

    \Lab_UT.didp.regrce1.q_esr_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20033\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22205\,
            ce => \N__12705\,
            sr => \N__20666\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__15494\,
            in2 => \N__17248\,
            in3 => \N__19865\,
            lcout => \Lab_UT.dictrl.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__19227\,
            in1 => \N__14978\,
            in2 => \N__14919\,
            in3 => \N__18628\,
            lcout => \Lab_UT.dictrl.G_25_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_4_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111111111"
        )
    port map (
            in0 => \N__18339\,
            in1 => \N__15774\,
            in2 => \N__12918\,
            in3 => \N__18441\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__19228\,
            in1 => \N__14724\,
            in2 => \N__12693\,
            in3 => \N__14979\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_25_i_a5_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100000101"
        )
    port map (
            in0 => \N__12729\,
            in1 => \N__18590\,
            in2 => \N__12690\,
            in3 => \N__15073\,
            lcout => \Lab_UT.un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19581\,
            in2 => \N__19256\,
            in3 => \N__19120\,
            lcout => \Lab_UT.dictrl.G_14_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19596\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18708\,
            in2 => \_gnd_net_\,
            in3 => \N__18338\,
            lcout => \Lab_UT.dictrl.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011111100"
        )
    port map (
            in0 => \N__15264\,
            in1 => \N__12744\,
            in2 => \N__12762\,
            in3 => \N__12939\,
            lcout => OPEN,
            ltout => \Lab_UT.i8_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_2_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12750\,
            in2 => \N__12765\,
            in3 => \N__18341\,
            lcout => \Lab_UT.didp.g0_0_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18550\,
            in1 => \N__21229\,
            in2 => \N__17247\,
            in3 => \N__19695\,
            lcout => \Lab_UT.dictrl.g0_0_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__19886\,
            in1 => \_gnd_net_\,
            in2 => \N__18469\,
            in3 => \N__20135\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__21481\,
            in1 => \N__19029\,
            in2 => \N__12753\,
            in3 => \N__21230\,
            lcout => \Lab_UT.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19600\,
            in1 => \N__17231\,
            in2 => \_gnd_net_\,
            in3 => \N__18549\,
            lcout => \Lab_UT.dictrl.g0_0_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__12738\,
            in1 => \N__14996\,
            in2 => \N__19281\,
            in3 => \N__12834\,
            lcout => \Lab_UT.dictrl.G_25_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19919\,
            in1 => \N__12723\,
            in2 => \N__12714\,
            in3 => \N__12924\,
            lcout => \Lab_UT.dictrl.N_57_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__20183\,
            in1 => \N__19400\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.m13_out\,
            ltout => \Lab_UT.dictrl.m13_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__21468\,
            in1 => \N__20152\,
            in2 => \N__12858\,
            in3 => \N__21212\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_18_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17243\,
            in1 => \N__12954\,
            in2 => \N__12855\,
            in3 => \N__19918\,
            lcout => \Lab_UT.dictrl.N_22_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19985\,
            in1 => \_gnd_net_\,
            in2 => \N__20157\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.g1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__17238\,
            in1 => \N__19607\,
            in2 => \N__18561\,
            in3 => \N__15681\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000001111"
        )
    port map (
            in0 => \N__12852\,
            in1 => \N__12846\,
            in2 => \N__12837\,
            in3 => \N__18348\,
            lcout => \Lab_UT.dictrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m34_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15398\,
            in2 => \_gnd_net_\,
            in3 => \N__19401\,
            lcout => \Lab_UT.dictrl.m34Z0Z_1\,
            ltout => \Lab_UT.dictrl.m34Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m34_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12810\,
            in1 => \N__13111\,
            in2 => \N__12828\,
            in3 => \N__15737\,
            lcout => \Lab_UT.dictrl.N_67_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_7_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15736\,
            in1 => \N__12809\,
            in2 => \N__13113\,
            in3 => \N__15589\,
            lcout => \Lab_UT.dictrl.g1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19740\,
            in2 => \_gnd_net_\,
            in3 => \N__19359\,
            lcout => \Lab_UT.dictrl.m22Z0Z_1\,
            ltout => \Lab_UT.dictrl.m22Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_8_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19989\,
            in1 => \N__15262\,
            in2 => \N__12957\,
            in3 => \N__21223\,
            lcout => \Lab_UT.dictrl.N_72_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15263\,
            in1 => \N__21104\,
            in2 => \N__12948\,
            in3 => \N__12938\,
            lcout => \Lab_UT.dictrl.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_4_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15665\,
            in1 => \N__15367\,
            in2 => \N__15645\,
            in3 => \N__15399\,
            lcout => \Lab_UT.dictrl.m22Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_8_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__15351\,
            in1 => \N__15320\,
            in2 => \N__15342\,
            in3 => \N__19921\,
            lcout => \Lab_UT.dictrl.g1_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__19739\,
            in1 => \N__19347\,
            in2 => \N__15439\,
            in3 => \N__15588\,
            lcout => \Lab_UT.dictrl.g0_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m5_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15400\,
            in1 => \N__13001\,
            in2 => \N__15376\,
            in3 => \N__15827\,
            lcout => \N_63_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_x1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15641\,
            in1 => \N__12899\,
            in2 => \N__12887\,
            in3 => \N__12869\,
            lcout => \Lab_UT.dictrl.g1_0_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_1_5_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15401\,
            in1 => \N__15815\,
            in2 => \N__12888\,
            in3 => \N__20192\,
            lcout => \Lab_UT.dictrl.g1_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__13002\,
            in1 => \_gnd_net_\,
            in2 => \N__15440\,
            in3 => \N__12870\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19348\,
            in1 => \N__15666\,
            in2 => \N__13125\,
            in3 => \N__13122\,
            lcout => \Lab_UT.dictrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_rep1_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13099\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22191\,
            ce => \N__20789\,
            sr => \N__20696\
        );

    \buart.Z_rx.shifter_7_rep1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13034\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22191\,
            ce => \N__20789\,
            sr => \N__20696\
        );

    \buart.Z_rx.shifter_fast_6_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22191\,
            ce => \N__20789\,
            sr => \N__20696\
        );

    \buart.Z_rx.shifter_fast_7_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22191\,
            ce => \N__20789\,
            sr => \N__20696\
        );

    \uu2.w_addr_displaying_fast_8_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110100"
        )
    port map (
            in0 => \N__12982\,
            in1 => \N__15878\,
            in2 => \N__16348\,
            in3 => \N__13422\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20627\
        );

    \uu2.w_addr_displaying_8_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000010"
        )
    port map (
            in0 => \N__15877\,
            in1 => \N__12981\,
            in2 => \N__13427\,
            in3 => \N__13242\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20627\
        );

    \uu2.w_addr_displaying_RNI0ES07_8_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011111111"
        )
    port map (
            in0 => \N__13241\,
            in1 => \N__13413\,
            in2 => \N__12990\,
            in3 => \N__21785\,
            lcout => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\,
            ltout => \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111101010000"
        )
    port map (
            in0 => \N__13417\,
            in1 => \_gnd_net_\,
            in2 => \N__12960\,
            in3 => \N__13372\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20627\
        );

    \uu2.w_addr_displaying_5_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__13373\,
            in1 => \N__15876\,
            in2 => \N__13305\,
            in3 => \N__13418\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20627\
        );

    \uu2.w_addr_displaying_ness_RNO_0_6_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__13295\,
            in1 => \_gnd_net_\,
            in2 => \N__13426\,
            in3 => \N__13371\,
            lcout => \uu2.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000011000"
        )
    port map (
            in0 => \N__13183\,
            in1 => \N__16603\,
            in2 => \N__13256\,
            in3 => \N__13293\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__13294\,
            in1 => \N__13240\,
            in2 => \N__16617\,
            in3 => \N__13184\,
            lcout => \uu2.bitmap_pmux_sn_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_290_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011101"
        )
    port map (
            in0 => \N__14657\,
            in1 => \N__14482\,
            in2 => \N__13468\,
            in3 => \N__13559\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \uu2.bitmap_194_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010101"
        )
    port map (
            in0 => \N__13558\,
            in1 => \N__13455\,
            in2 => \N__14491\,
            in3 => \N__14656\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \uu2.bitmap_66_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__14659\,
            in1 => \N__14486\,
            in2 => \N__13469\,
            in3 => \N__13561\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \uu2.bitmap_RNIPDM31_66_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__13149\,
            in1 => \N__16602\,
            in2 => \N__16541\,
            in3 => \N__13143\,
            lcout => \uu2.bitmap_pmux_20_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__14655\,
            in1 => \N__14478\,
            in2 => \N__13467\,
            in3 => \N__13557\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \uu2.bitmap_34_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__13560\,
            in1 => \N__13459\,
            in2 => \N__14492\,
            in3 => \N__14658\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \uu2.bitmap_RNIP2JO1_34_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111010"
        )
    port map (
            in0 => \N__13803\,
            in1 => \N__13797\,
            in2 => \N__13791\,
            in3 => \N__13749\,
            lcout => \uu2.bitmap_RNIP2JO1Z0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_69_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__13562\,
            in1 => \N__13463\,
            in2 => \N__14493\,
            in3 => \N__14660\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20625\
        );

    \Lab_UT.dictrl.next_state_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011000000"
        )
    port map (
            in0 => \N__14787\,
            in1 => \N__18480\,
            in2 => \N__14760\,
            in3 => \N__18347\,
            lcout => \Lab_UT.dictrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22256\,
            ce => \N__18771\,
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17797\,
            in1 => \N__13728\,
            in2 => \_gnd_net_\,
            in3 => \N__13682\,
            lcout => \Lab_UT.sec2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13649\,
            in1 => \N__14360\,
            in2 => \_gnd_net_\,
            in3 => \N__17798\,
            lcout => \Lab_UT.sec2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__16697\,
            in2 => \_gnd_net_\,
            in3 => \N__13620\,
            lcout => \Lab_UT.min2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13590\,
            in1 => \N__17100\,
            in2 => \_gnd_net_\,
            in3 => \N__17800\,
            lcout => \Lab_UT.min1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13536\,
            in1 => \N__13509\,
            in2 => \_gnd_net_\,
            in3 => \N__17799\,
            lcout => \Lab_UT.min1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__13827\,
            in1 => \N__14372\,
            in2 => \N__14115\,
            in3 => \N__14064\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \uu2.bitmap_RNIOPSS_212_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__14037\,
            in1 => \N__16405\,
            in2 => \N__14019\,
            in3 => \N__14031\,
            lcout => \uu2.bitmap_pmux_17_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_0_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15880\,
            in2 => \_gnd_net_\,
            in3 => \N__14017\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \uu2.bitmap_RNI65TM_72_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__13983\,
            in1 => \N__16404\,
            in2 => \N__14018\,
            in3 => \N__13989\,
            lcout => \uu2.bitmap_pmux_16_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_7_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__16406\,
            in1 => \N__15881\,
            in2 => \_gnd_net_\,
            in3 => \N__15917\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \uu2.bitmap_72_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__13964\,
            in1 => \N__13936\,
            in2 => \N__14150\,
            in3 => \N__13898\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \uu2.bitmap_200_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__13896\,
            in1 => \N__14133\,
            in2 => \N__13945\,
            in3 => \N__13962\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \uu2.bitmap_296_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__13963\,
            in1 => \N__13935\,
            in2 => \N__14149\,
            in3 => \N__13897\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20622\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17796\,
            in1 => \N__13872\,
            in2 => \_gnd_net_\,
            in3 => \N__14591\,
            lcout => \Lab_UT.sec1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14520\,
            in1 => \N__17025\,
            in2 => \_gnd_net_\,
            in3 => \N__17795\,
            lcout => \Lab_UT.min1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17794\,
            in1 => \N__14451\,
            in2 => \_gnd_net_\,
            in3 => \N__14421\,
            lcout => \Lab_UT.sec1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_2_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14356\,
            in2 => \_gnd_net_\,
            in3 => \N__17892\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__14301\,
            in1 => \N__20932\,
            in2 => \N__14262\,
            in3 => \N__16983\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__16984\,
            in1 => \N__14242\,
            in2 => \N__14217\,
            in3 => \N__14214\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16880\,
            in1 => \N__17300\,
            in2 => \N__16706\,
            in3 => \N__16748\,
            lcout => \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__16878\,
            in1 => \N__14681\,
            in2 => \N__17611\,
            in3 => \N__14602\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14603\,
            in1 => \N__17786\,
            in2 => \_gnd_net_\,
            in3 => \N__16879\,
            lcout => \Lab_UT.min2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17603\,
            in1 => \_gnd_net_\,
            in2 => \N__17802\,
            in3 => \N__14682\,
            lcout => \Lab_UT.min1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21389\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22233\,
            ce => \N__14628\,
            sr => \N__20672\
        );

    \Lab_UT.dispString.dOut_RNO_3_1_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18206\,
            in1 => \N__18092\,
            in2 => \N__17998\,
            in3 => \N__14604\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110000"
        )
    port map (
            in0 => \N__14592\,
            in1 => \N__18093\,
            in2 => \N__14562\,
            in3 => \N__14533\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18202\,
            lcout => \Lab_UT.dispString.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19507\,
            in1 => \N__19883\,
            in2 => \N__18468\,
            in3 => \N__18330\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20750\,
            lcout => \Lab_UT.bu_rx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__15074\,
            in1 => \N__15027\,
            in2 => \N__14826\,
            in3 => \N__14998\,
            lcout => \Lab_UT.dictrl.dicLdAMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22227\,
            ce => 'H',
            sr => \N__20670\
        );

    \Lab_UT.dictrl.state_ret_5_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__14999\,
            in1 => \N__15075\,
            in2 => \N__18363\,
            in3 => \N__18592\,
            lcout => \Lab_UT.dictrl.dicRun_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22227\,
            ce => 'H',
            sr => \N__20670\
        );

    \Lab_UT.dictrl.state_ret_9_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__18591\,
            in1 => \N__15028\,
            in2 => \N__19133\,
            in3 => \N__15000\,
            lcout => \Lab_UT.dicLdSones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22227\,
            ce => 'H',
            sr => \N__20670\
        );

    \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18445\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__14822\,
            lcout => \Lab_UT.LdAMones\,
            ltout => \Lab_UT.LdAMones_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14843\,
            in1 => \N__18239\,
            in2 => \N__14799\,
            in3 => \N__14850\,
            lcout => \Lab_UT.loadalarm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__14690\,
            in1 => \N__15308\,
            in2 => \_gnd_net_\,
            in3 => \N__14796\,
            lcout => \Lab_UT.next_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI81O17_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__19282\,
            in1 => \N__15773\,
            in2 => \N__14720\,
            in3 => \N__18421\,
            lcout => \Lab_UT.dictrl.g0_1_mb_rn_0\,
            ltout => \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__14691\,
            in1 => \_gnd_net_\,
            in2 => \N__14790\,
            in3 => \N__15309\,
            lcout => \Lab_UT.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22220\,
            ce => \N__18507\,
            sr => \N__20663\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__18299\,
            in1 => \N__14783\,
            in2 => \N__14753\,
            in3 => \N__18423\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14716\,
            in2 => \N__14694\,
            in3 => \N__19286\,
            lcout => \Lab_UT.dictrl.state_i_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22220\,
            ce => \N__18507\,
            sr => \N__20663\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__18298\,
            in1 => \_gnd_net_\,
            in2 => \N__19293\,
            in3 => \N__18422\,
            lcout => \Lab_UT.dictrl.g0_1_mb_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18700\,
            in2 => \_gnd_net_\,
            in3 => \N__18297\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un15_loadalarm_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__19103\,
            in1 => \N__18420\,
            in2 => \N__14853\,
            in3 => \N__19459\,
            lcout => \Lab_UT.dictrl.loadalarm_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18930\,
            in1 => \N__17907\,
            in2 => \N__18824\,
            in3 => \N__15195\,
            lcout => \Lab_UT.next_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15198\,
            in1 => \N__18823\,
            in2 => \N__18939\,
            in3 => \N__17910\,
            lcout => \Lab_UT.dictrl.state_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18931\,
            in1 => \N__17908\,
            in2 => \N__18825\,
            in3 => \N__15196\,
            lcout => \Lab_UT.dictrl.state_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15197\,
            in1 => \N__18822\,
            in2 => \N__18938\,
            in3 => \N__17909\,
            lcout => \Lab_UT.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18419\,
            in1 => \N__19458\,
            in2 => \N__15111\,
            in3 => \N__19831\,
            lcout => \Lab_UT.LdAStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__18671\,
            in1 => \_gnd_net_\,
            in2 => \N__18654\,
            in3 => \N__19254\,
            lcout => \Lab_UT.state_i_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19253\,
            in1 => \N__18650\,
            in2 => \_gnd_net_\,
            in3 => \N__18670\,
            lcout => \Lab_UT.dictrl.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__17164\,
            in1 => \N__17141\,
            in2 => \N__19628\,
            in3 => \N__19255\,
            lcout => \Lab_UT_dictrl_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => \N__18515\,
            sr => \N__20671\
        );

    \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__19247\,
            in1 => \N__15152\,
            in2 => \N__15138\,
            in3 => \N__15112\,
            lcout => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__15114\,
            in1 => \N__19595\,
            in2 => \N__17168\,
            in3 => \N__15153\,
            lcout => \Lab_UT.dictrl.next_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22206\,
            ce => \N__18748\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__14870\,
            in1 => \N__15164\,
            in2 => \N__15126\,
            in3 => \N__19471\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_20_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__15113\,
            in1 => \N__19593\,
            in2 => \N__15090\,
            in3 => \N__15087\,
            lcout => OPEN,
            ltout => \Lab_UT.next_state_1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__15063\,
            in1 => \N__14877\,
            in2 => \N__15036\,
            in3 => \N__15033\,
            lcout => \Lab_UT.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14980\,
            in1 => \N__14925\,
            in2 => \N__14915\,
            in3 => \N__19248\,
            lcout => \Lab_UT.didp.g0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__14871\,
            in1 => \N__15165\,
            in2 => \N__19508\,
            in3 => \N__18684\,
            lcout => \Lab_UT.dictrl.N_20\,
            ltout => \Lab_UT.dictrl.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__19252\,
            in1 => \N__19594\,
            in2 => \N__14856\,
            in3 => \N__17140\,
            lcout => \Lab_UT.next_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18455\,
            in2 => \_gnd_net_\,
            in3 => \N__19888\,
            lcout => \Lab_UT.dictrl.m34_0\,
            ltout => \Lab_UT.dictrl.m34_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m35_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__15281\,
            in1 => \N__15490\,
            in2 => \N__15231\,
            in3 => \N__18336\,
            lcout => \Lab_UT.dictrl.next_state_1_3\,
            ltout => \Lab_UT.dictrl.next_state_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__18629\,
            in1 => \_gnd_net_\,
            in2 => \N__15228\,
            in3 => \N__19231\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19229\,
            in1 => \N__19601\,
            in2 => \_gnd_net_\,
            in3 => \N__18334\,
            lcout => \Lab_UT.dictrl.N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__18335\,
            in1 => \N__19230\,
            in2 => \N__19622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__19887\,
            in1 => \N__15171\,
            in2 => \N__15201\,
            in3 => \N__15288\,
            lcout => \Lab_UT.dictrl.N_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__18337\,
            in1 => \N__15180\,
            in2 => \N__15495\,
            in3 => \N__15282\,
            lcout => \Lab_UT.dictrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22200\,
            ce => \N__18764\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__21466\,
            in1 => \N__15456\,
            in2 => \N__20140\,
            in3 => \N__18901\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19027\,
            in1 => \N__15273\,
            in2 => \N__15174\,
            in3 => \N__18902\,
            lcout => \Lab_UT.dictrl.N_60_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001100110"
        )
    port map (
            in0 => \N__19920\,
            in1 => \N__20058\,
            in2 => \N__15486\,
            in3 => \N__18345\,
            lcout => \Lab_UT.dictrl.m19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__15457\,
            in1 => \N__21095\,
            in2 => \_gnd_net_\,
            in3 => \N__21467\,
            lcout => OPEN,
            ltout => \N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001000"
        )
    port map (
            in0 => \N__19605\,
            in1 => \N__19134\,
            in2 => \N__15294\,
            in3 => \N__19496\,
            lcout => \Lab_UT.dictrl.G_6_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__21465\,
            in2 => \N__18913\,
            in3 => \N__18981\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__15237\,
            in1 => \N__19028\,
            in2 => \N__15291\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_59_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__18557\,
            in1 => \N__19606\,
            in2 => \N__17253\,
            in3 => \N__18982\,
            lcout => \Lab_UT.dictrl.i8_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111101"
        )
    port map (
            in0 => \N__21437\,
            in1 => \N__15458\,
            in2 => \N__18905\,
            in3 => \N__20127\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_x1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19338\,
            in1 => \N__21214\,
            in2 => \N__19775\,
            in3 => \N__19687\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m22_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_ns_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15267\,
            in3 => \N__15258\,
            lcout => \Lab_UT.dictrl.N_72_mux\,
            ltout => \Lab_UT.dictrl.N_72_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20125\,
            in2 => \N__15240\,
            in3 => \N__21436\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m7_a0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20196\,
            in2 => \_gnd_net_\,
            in3 => \N__19391\,
            lcout => m7_a0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__19392\,
            in1 => \N__18887\,
            in2 => \N__20204\,
            in3 => \N__20126\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__21435\,
            in1 => \_gnd_net_\,
            in2 => \N__15498\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m7_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21438\,
            lcout => \Lab_UT.dictrl.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_4_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15643\,
            in1 => \N__15668\,
            in2 => \N__18904\,
            in3 => \N__15377\,
            lcout => \Lab_UT.dictrl.g0_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__18886\,
            in1 => \N__19756\,
            in2 => \_gnd_net_\,
            in3 => \N__19345\,
            lcout => \Lab_UT.dictrl.gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15642\,
            in1 => \N__15667\,
            in2 => \N__15441\,
            in3 => \N__15408\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__15378\,
            in1 => \_gnd_net_\,
            in2 => \N__15354\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.g0_6_3\,
            ltout => \Lab_UT.dictrl.g0_6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19885\,
            in1 => \N__15341\,
            in2 => \N__15327\,
            in3 => \N__15324\,
            lcout => \Lab_UT.dictrl.N_57_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17184\,
            in1 => \N__15831\,
            in2 => \N__15816\,
            in3 => \N__20205\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15798\,
            in3 => \N__15795\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15789\,
            in1 => \N__15783\,
            in2 => \N__15777\,
            in3 => \N__19884\,
            lcout => \Lab_UT.dictrl.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19773\,
            in1 => \N__19698\,
            in2 => \N__18903\,
            in3 => \N__15611\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_10_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15618\,
            in1 => \N__19346\,
            in2 => \N__15750\,
            in3 => \N__15740\,
            lcout => \Lab_UT.dictrl.N_72_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_11_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15669\,
            in2 => \_gnd_net_\,
            in3 => \N__15644\,
            lcout => \Lab_UT.dictrl.g0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_rep1_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15612\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22194\,
            ce => \N__20791\,
            sr => \N__20697\
        );

    \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16134\,
            in1 => \N__20333\,
            in2 => \N__15528\,
            in3 => \N__16232\,
            lcout => \uu2.un3_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16234\,
            in1 => \N__16139\,
            in2 => \N__20342\,
            in3 => \N__21839\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15960\,
            sr => \N__15948\
        );

    \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15973\,
            in1 => \N__16153\,
            in2 => \_gnd_net_\,
            in3 => \N__21837\,
            lcout => OPEN,
            ltout => \uu2.un3_w_addr_user_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIINVH_4_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16192\,
            in1 => \N__16299\,
            in2 => \N__16269\,
            in3 => \N__16266\,
            lcout => \uu2.un3_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20340\,
            in1 => \N__21838\,
            in2 => \N__16140\,
            in3 => \N__16233\,
            lcout => \uu2.un404_ci\,
            ltout => \uu2.un404_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_7_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16154\,
            in1 => \N__16040\,
            in2 => \N__16197\,
            in3 => \N__16194\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15960\,
            sr => \N__15948\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16135\,
            in1 => \N__21786\,
            in2 => \_gnd_net_\,
            in3 => \N__16122\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__16041\,
            in1 => \N__16001\,
            in2 => \N__15990\,
            in3 => \N__15974\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15960\,
            sr => \N__15948\
        );

    \uu2.w_addr_displaying_7_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__15867\,
            in1 => \N__15918\,
            in2 => \_gnd_net_\,
            in3 => \N__16616\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20628\
        );

    \uu2.w_addr_displaying_0_rep1_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15866\,
            in2 => \_gnd_net_\,
            in3 => \N__16529\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20628\
        );

    \uu2.bitmap_111_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17547\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20628\
        );

    \uu2.bitmap_314_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011101"
        )
    port map (
            in0 => \N__16911\,
            in1 => \N__17708\,
            in2 => \N__16446\,
            in3 => \N__16473\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20626\
        );

    \uu2.bitmap_218_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010101"
        )
    port map (
            in0 => \N__16472\,
            in1 => \N__16432\,
            in2 => \N__17718\,
            in3 => \N__16910\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20626\
        );

    \uu2.bitmap_90_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__16913\,
            in1 => \N__17712\,
            in2 => \N__16447\,
            in3 => \N__16475\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20626\
        );

    \uu2.bitmap_RNIJ4K41_90_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__16601\,
            in1 => \N__16563\,
            in2 => \N__16540\,
            in3 => \N__16497\,
            lcout => \uu2.bitmap_pmux_19_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__16909\,
            in1 => \N__17704\,
            in2 => \N__16445\,
            in3 => \N__16471\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20626\
        );

    \uu2.bitmap_58_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__16474\,
            in1 => \N__16436\,
            in2 => \N__17719\,
            in3 => \N__16912\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20626\
        );

    \uu2.bitmap_RNIKGSI_58_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16403\,
            in1 => \N__16383\,
            in2 => \_gnd_net_\,
            in3 => \N__16377\,
            lcout => OPEN,
            ltout => \uu2.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIM5E21_314_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16370\,
            in2 => \N__16356\,
            in3 => \N__16347\,
            lcout => \uu2.bitmap_RNIM5E21Z0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__16662\,
            in1 => \N__16668\,
            in2 => \N__17370\,
            in3 => \N__16702\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16882\,
            in2 => \_gnd_net_\,
            in3 => \N__17299\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17329\,
            in1 => \N__20933\,
            in2 => \N__16764\,
            in3 => \N__16742\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__16743\,
            in1 => \N__17359\,
            in2 => \N__16761\,
            in3 => \N__16661\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17028\,
            in2 => \_gnd_net_\,
            in3 => \N__17102\,
            lcout => \Lab_UT.didp.reset_12_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16741\,
            in1 => \N__16881\,
            in2 => \_gnd_net_\,
            in3 => \N__17298\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17328\,
            in1 => \N__21134\,
            in2 => \N__16710\,
            in3 => \N__16701\,
            lcout => \Lab_UT.didp.countrce3.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNIBN0Q1_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17399\,
            in2 => \_gnd_net_\,
            in3 => \N__17330\,
            lcout => \Lab_UT.didp.un1_dicLdMones_0\,
            ltout => \Lab_UT.didp.un1_dicLdMones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__16883\,
            in1 => \N__16851\,
            in2 => \N__16650\,
            in3 => \N__17358\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0_sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__17316\,
            in1 => \N__20051\,
            in2 => \_gnd_net_\,
            in3 => \N__17292\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIFV4E_1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18112\,
            in2 => \_gnd_net_\,
            in3 => \N__18207\,
            lcout => \Lab_UT.dispString.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__21395\,
            in1 => \N__17026\,
            in2 => \N__17676\,
            in3 => \N__17103\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17027\,
            in1 => \N__16838\,
            in2 => \N__17040\,
            in3 => \N__16781\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16978\,
            in1 => \N__17773\,
            in2 => \_gnd_net_\,
            in3 => \N__16947\,
            lcout => \Lab_UT.sec2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__17293\,
            in1 => \N__16884\,
            in2 => \N__21396\,
            in3 => \N__17317\,
            lcout => \Lab_UT.didp.countrce3.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__16780\,
            in1 => \N__17610\,
            in2 => \N__17580\,
            in3 => \N__16842\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNIHGGI1_3_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16809\,
            in2 => \_gnd_net_\,
            in3 => \N__17675\,
            lcout => \Lab_UT.didp.un1_dicLdMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17882\,
            in1 => \N__17832\,
            in2 => \_gnd_net_\,
            in3 => \N__17774\,
            lcout => \Lab_UT.sec2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17674\,
            in1 => \N__20926\,
            in2 => \N__17631\,
            in3 => \N__17609\,
            lcout => \Lab_UT.didp.countrce4.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17558\,
            in2 => \_gnd_net_\,
            in3 => \N__17535\,
            lcout => \oneSecStrb\,
            ltout => \oneSecStrb_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIKUO21_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001001"
        )
    port map (
            in0 => \N__18117\,
            in1 => \N__17980\,
            in2 => \N__17433\,
            in3 => \N__18222\,
            lcout => \Lab_UT.dispString.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001001"
        )
    port map (
            in0 => \N__17403\,
            in1 => \N__17376\,
            in2 => \N__17369\,
            in3 => \N__17331\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000110111"
        )
    port map (
            in0 => \N__19287\,
            in1 => \N__19148\,
            in2 => \N__18804\,
            in3 => \N__19055\,
            lcout => \Lab_UT.dictrl.state_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22228\,
            ce => \N__18519\,
            sr => \N__20667\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100011101"
        )
    port map (
            in0 => \N__19056\,
            in1 => \N__18803\,
            in2 => \N__19152\,
            in3 => \N__19288\,
            lcout => \Lab_UT.dictrl.state_ret_2_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22228\,
            ce => \N__18519\,
            sr => \N__20667\
        );

    \Lab_UT.dictrl.state_ret_6_ess_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000111111101"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__19289\,
            in2 => \N__19629\,
            in3 => \N__17145\,
            lcout => \Lab_UT.dictrl.state_i_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22228\,
            ce => \N__18519\,
            sr => \N__20667\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18704\,
            in2 => \_gnd_net_\,
            in3 => \N__18301\,
            lcout => \Lab_UT.dictrl.m19_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_esr_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19290\,
            in1 => \N__18672\,
            in2 => \N__18649\,
            in3 => \N__18602\,
            lcout => \Lab_UT.dictrl.next_state66_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22228\,
            ce => \N__18519\,
            sr => \N__20667\
        );

    \Lab_UT.dictrl.state_ret_5_RNICG571_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18418\,
            in1 => \N__18359\,
            in2 => \_gnd_net_\,
            in3 => \N__18300\,
            lcout => \Lab_UT.LdASones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__17975\,
            in1 => \N__18221\,
            in2 => \_gnd_net_\,
            in3 => \N__18118\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__20673\
        );

    \Lab_UT.dictrl.g1_8_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19776\,
            in1 => \N__19361\,
            in2 => \N__18914\,
            in3 => \N__19697\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20095\,
            in1 => \N__17928\,
            in2 => \N__17916\,
            in3 => \N__19864\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_14_0_a2_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__19257\,
            in2 => \N__17913\,
            in3 => \N__18950\,
            lcout => \Lab_UT.dictrl.G_14_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__19360\,
            in1 => \N__18906\,
            in2 => \_gnd_net_\,
            in3 => \N__19777\,
            lcout => OPEN,
            ltout => \shifter_1_rep1_RNI0FPF_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__19863\,
            in1 => \N__20094\,
            in2 => \N__18954\,
            in3 => \N__21494\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__18951\,
            in1 => \N__21152\,
            in2 => \N__18942\,
            in3 => \N__19460\,
            lcout => \Lab_UT.dictrl.G_14_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__19778\,
            in1 => \N__21495\,
            in2 => \N__18915\,
            in3 => \N__19362\,
            lcout => OPEN,
            ltout => \N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100010"
        )
    port map (
            in0 => \N__18837\,
            in1 => \N__21153\,
            in2 => \N__18828\,
            in3 => \N__19461\,
            lcout => \Lab_UT.dictrl.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__19618\,
            in1 => \N__20214\,
            in2 => \N__19164\,
            in3 => \N__19136\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18799\,
            in1 => \_gnd_net_\,
            in2 => \N__18774\,
            in3 => \N__18714\,
            lcout => \Lab_UT.dictrl.next_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22207\,
            ce => \N__18763\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m14_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__21091\,
            in1 => \N__21492\,
            in2 => \_gnd_net_\,
            in3 => \N__19041\,
            lcout => \Lab_UT.dictrl.N_15_0\,
            ltout => \Lab_UT.dictrl.N_15_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111011"
        )
    port map (
            in0 => \N__21093\,
            in1 => \N__20229\,
            in2 => \N__18720\,
            in3 => \N__19506\,
            lcout => \Lab_UT.dictrl.N_60\,
            ltout => \Lab_UT.dictrl.N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18962\,
            in2 => \N__18717\,
            in3 => \N__19917\,
            lcout => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__19305\,
            in1 => \N__19291\,
            in2 => \_gnd_net_\,
            in3 => \N__19916\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__18963\,
            in1 => \N__19292\,
            in2 => \N__19167\,
            in3 => \N__19163\,
            lcout => \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101110000"
        )
    port map (
            in0 => \N__19500\,
            in1 => \N__19135\,
            in2 => \N__19627\,
            in3 => \N__19910\,
            lcout => \Lab_UT.dictrl.G_6_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__21237\,
            in1 => \N__20874\,
            in2 => \N__21379\,
            in3 => \N__21486\,
            lcout => OPEN,
            ltout => \G_6_0_a6_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001000100"
        )
    port map (
            in0 => \N__18999\,
            in1 => \N__19617\,
            in2 => \N__19077\,
            in3 => \N__19074\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19407\,
            in2 => \N__19068\,
            in3 => \N__19065\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_5_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110011011"
        )
    port map (
            in0 => \N__19909\,
            in1 => \N__21236\,
            in2 => \N__21493\,
            in3 => \N__19040\,
            lcout => \Lab_UT.dictrl.next_state_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__19501\,
            in1 => \N__18998\,
            in2 => \_gnd_net_\,
            in3 => \N__18986\,
            lcout => \Lab_UT.dictrl.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__19935\,
            in1 => \N__20228\,
            in2 => \N__21135\,
            in3 => \N__19502\,
            lcout => \Lab_UT.dictrl.i8_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__21234\,
            in1 => \N__20203\,
            in2 => \N__20156\,
            in3 => \N__19393\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20061\,
            in3 => \N__21482\,
            lcout => \Lab_UT.dictrl.N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_4_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20007\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_3_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101010101"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__19640\,
            in2 => \N__19944\,
            in3 => \N__19941\,
            lcout => \Lab_UT.dictrl.i9_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19927\,
            in1 => \N__21235\,
            in2 => \N__19779\,
            in3 => \N__19691\,
            lcout => OPEN,
            ltout => \G_6_0_a6_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__19641\,
            in1 => \N__19626\,
            in2 => \N__19515\,
            in3 => \N__19512\,
            lcout => \Lab_UT.dictrl.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20848\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__20796\,
            sr => \N__20698\
        );

    \buart.Z_rx.shifter_1_rep1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__20796\,
            sr => \N__20698\
        );

    \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__20846\,
            in1 => \N__21480\,
            in2 => \N__21335\,
            in3 => \N__21233\,
            lcout => \N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21115\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__20796\,
            sr => \N__20698\
        );

    \buart.Z_tx.bitcount_1_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111111100"
        )
    port map (
            in0 => \N__21522\,
            in1 => \N__21558\,
            in2 => \N__20463\,
            in3 => \N__21583\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => 'H',
            sr => \N__20699\
        );

    \buart.Z_tx.bitcount_0_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21581\,
            in1 => \N__20461\,
            in2 => \_gnd_net_\,
            in3 => \N__21521\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => 'H',
            sr => \N__20699\
        );

    \buart.Z_tx.bitcount_3_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__21603\,
            in1 => \N__21501\,
            in2 => \N__21588\,
            in3 => \N__20457\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => 'H',
            sr => \N__20699\
        );

    \buart.Z_tx.bitcount_2_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100100000110"
        )
    port map (
            in0 => \N__21582\,
            in1 => \N__21609\,
            in2 => \N__20462\,
            in3 => \N__21540\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => 'H',
            sr => \N__20699\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20453\,
            in2 => \_gnd_net_\,
            in3 => \N__21580\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20343\,
            in1 => \N__21805\,
            in2 => \_gnd_net_\,
            in3 => \N__20301\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21807\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21879\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21840\,
            in1 => \N__21806\,
            in2 => \_gnd_net_\,
            in3 => \N__21693\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__21519\,
            in1 => \N__21556\,
            in2 => \_gnd_net_\,
            in3 => \N__21584\,
            lcout => \buart.Z_tx.un1_bitcount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21954\,
            in2 => \_gnd_net_\,
            in3 => \N__21938\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21937\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21602\,
            in2 => \_gnd_net_\,
            in3 => \N__21518\,
            lcout => OPEN,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__21538\,
            in1 => \N__21555\,
            in2 => \N__21591\,
            in3 => \N__21894\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__21557\,
            in1 => \N__21539\,
            in2 => \N__21525\,
            in3 => \N__21520\,
            lcout => \buart.Z_tx.un1_bitcount_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21953\,
            in2 => \N__21939\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21918\,
            in3 => \N__22296\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__22274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21896\,
            in1 => \N__21963\,
            in2 => \_gnd_net_\,
            in3 => \N__22293\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__22274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21990\,
            in3 => \N__22290\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__22274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__21897\,
            in1 => \_gnd_net_\,
            in2 => \N__22002\,
            in3 => \N__22287\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__22274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21977\,
            in1 => \N__21895\,
            in2 => \_gnd_net_\,
            in3 => \N__22284\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__21986\,
            in2 => \N__21978\,
            in3 => \N__21962\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21952\,
            in1 => \N__21933\,
            in2 => \N__21917\,
            in3 => \N__21903\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
