// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 19 2019 07:10:59

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__19573;
    wire N__19572;
    wire N__19571;
    wire N__19564;
    wire N__19563;
    wire N__19562;
    wire N__19555;
    wire N__19554;
    wire N__19553;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19537;
    wire N__19536;
    wire N__19535;
    wire N__19528;
    wire N__19527;
    wire N__19526;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19501;
    wire N__19500;
    wire N__19499;
    wire N__19492;
    wire N__19491;
    wire N__19490;
    wire N__19473;
    wire N__19472;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19451;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19436;
    wire N__19435;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19429;
    wire N__19428;
    wire N__19425;
    wire N__19424;
    wire N__19423;
    wire N__19422;
    wire N__19417;
    wire N__19414;
    wire N__19407;
    wire N__19400;
    wire N__19397;
    wire N__19390;
    wire N__19387;
    wire N__19382;
    wire N__19371;
    wire N__19368;
    wire N__19367;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19351;
    wire N__19350;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19335;
    wire N__19330;
    wire N__19329;
    wire N__19324;
    wire N__19319;
    wire N__19314;
    wire N__19313;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19301;
    wire N__19296;
    wire N__19287;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19282;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19265;
    wire N__19264;
    wire N__19261;
    wire N__19260;
    wire N__19257;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19203;
    wire N__19198;
    wire N__19195;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19174;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19147;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19137;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19104;
    wire N__19099;
    wire N__19096;
    wire N__19091;
    wire N__19088;
    wire N__19083;
    wire N__19074;
    wire N__19073;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19069;
    wire N__19068;
    wire N__19065;
    wire N__19060;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19048;
    wire N__19045;
    wire N__19040;
    wire N__19039;
    wire N__19038;
    wire N__19037;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19025;
    wire N__19024;
    wire N__19021;
    wire N__19014;
    wire N__19011;
    wire N__19006;
    wire N__19001;
    wire N__18998;
    wire N__18987;
    wire N__18984;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18972;
    wire N__18969;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18960;
    wire N__18959;
    wire N__18956;
    wire N__18955;
    wire N__18954;
    wire N__18953;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18938;
    wire N__18933;
    wire N__18928;
    wire N__18925;
    wire N__18918;
    wire N__18909;
    wire N__18908;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18902;
    wire N__18901;
    wire N__18900;
    wire N__18897;
    wire N__18896;
    wire N__18895;
    wire N__18894;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18878;
    wire N__18877;
    wire N__18874;
    wire N__18865;
    wire N__18858;
    wire N__18855;
    wire N__18846;
    wire N__18845;
    wire N__18844;
    wire N__18843;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18798;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18777;
    wire N__18776;
    wire N__18775;
    wire N__18772;
    wire N__18767;
    wire N__18766;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18747;
    wire N__18746;
    wire N__18745;
    wire N__18744;
    wire N__18743;
    wire N__18742;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18719;
    wire N__18714;
    wire N__18713;
    wire N__18712;
    wire N__18711;
    wire N__18710;
    wire N__18709;
    wire N__18708;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18704;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18700;
    wire N__18699;
    wire N__18698;
    wire N__18697;
    wire N__18696;
    wire N__18695;
    wire N__18694;
    wire N__18693;
    wire N__18692;
    wire N__18691;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18668;
    wire N__18667;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18663;
    wire N__18662;
    wire N__18661;
    wire N__18660;
    wire N__18659;
    wire N__18658;
    wire N__18657;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18653;
    wire N__18652;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18648;
    wire N__18645;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18527;
    wire N__18526;
    wire N__18523;
    wire N__18522;
    wire N__18517;
    wire N__18512;
    wire N__18507;
    wire N__18506;
    wire N__18505;
    wire N__18504;
    wire N__18503;
    wire N__18502;
    wire N__18501;
    wire N__18500;
    wire N__18499;
    wire N__18498;
    wire N__18497;
    wire N__18496;
    wire N__18495;
    wire N__18494;
    wire N__18493;
    wire N__18492;
    wire N__18491;
    wire N__18490;
    wire N__18489;
    wire N__18488;
    wire N__18487;
    wire N__18486;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18481;
    wire N__18480;
    wire N__18479;
    wire N__18478;
    wire N__18477;
    wire N__18476;
    wire N__18475;
    wire N__18474;
    wire N__18473;
    wire N__18472;
    wire N__18471;
    wire N__18470;
    wire N__18469;
    wire N__18468;
    wire N__18467;
    wire N__18466;
    wire N__18465;
    wire N__18464;
    wire N__18463;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18459;
    wire N__18458;
    wire N__18457;
    wire N__18456;
    wire N__18455;
    wire N__18454;
    wire N__18453;
    wire N__18452;
    wire N__18451;
    wire N__18450;
    wire N__18449;
    wire N__18448;
    wire N__18447;
    wire N__18446;
    wire N__18445;
    wire N__18444;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18440;
    wire N__18439;
    wire N__18438;
    wire N__18437;
    wire N__18436;
    wire N__18435;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18426;
    wire N__18425;
    wire N__18424;
    wire N__18423;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18235;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18206;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18171;
    wire N__18170;
    wire N__18167;
    wire N__18166;
    wire N__18163;
    wire N__18162;
    wire N__18161;
    wire N__18160;
    wire N__18159;
    wire N__18158;
    wire N__18157;
    wire N__18150;
    wire N__18145;
    wire N__18142;
    wire N__18137;
    wire N__18130;
    wire N__18127;
    wire N__18122;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18095;
    wire N__18092;
    wire N__18091;
    wire N__18090;
    wire N__18089;
    wire N__18088;
    wire N__18087;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18069;
    wire N__18062;
    wire N__18055;
    wire N__18046;
    wire N__18037;
    wire N__18030;
    wire N__18027;
    wire N__18026;
    wire N__18025;
    wire N__18022;
    wire N__18021;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18015;
    wire N__18012;
    wire N__18007;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17986;
    wire N__17981;
    wire N__17974;
    wire N__17971;
    wire N__17966;
    wire N__17961;
    wire N__17958;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17946;
    wire N__17945;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17928;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17895;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17887;
    wire N__17886;
    wire N__17881;
    wire N__17878;
    wire N__17877;
    wire N__17876;
    wire N__17875;
    wire N__17874;
    wire N__17871;
    wire N__17870;
    wire N__17865;
    wire N__17862;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17856;
    wire N__17849;
    wire N__17846;
    wire N__17841;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17765;
    wire N__17760;
    wire N__17757;
    wire N__17756;
    wire N__17753;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17742;
    wire N__17741;
    wire N__17740;
    wire N__17739;
    wire N__17736;
    wire N__17731;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17704;
    wire N__17703;
    wire N__17702;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17687;
    wire N__17686;
    wire N__17683;
    wire N__17674;
    wire N__17669;
    wire N__17664;
    wire N__17661;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17616;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17547;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17529;
    wire N__17526;
    wire N__17525;
    wire N__17522;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17454;
    wire N__17453;
    wire N__17452;
    wire N__17451;
    wire N__17450;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17425;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17411;
    wire N__17410;
    wire N__17409;
    wire N__17406;
    wire N__17405;
    wire N__17404;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17376;
    wire N__17373;
    wire N__17372;
    wire N__17369;
    wire N__17368;
    wire N__17367;
    wire N__17366;
    wire N__17361;
    wire N__17358;
    wire N__17353;
    wire N__17350;
    wire N__17345;
    wire N__17340;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17326;
    wire N__17323;
    wire N__17318;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17274;
    wire N__17273;
    wire N__17270;
    wire N__17269;
    wire N__17268;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17242;
    wire N__17235;
    wire N__17234;
    wire N__17231;
    wire N__17230;
    wire N__17229;
    wire N__17228;
    wire N__17227;
    wire N__17224;
    wire N__17219;
    wire N__17214;
    wire N__17211;
    wire N__17204;
    wire N__17199;
    wire N__17198;
    wire N__17197;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17186;
    wire N__17183;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17168;
    wire N__17165;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17127;
    wire N__17124;
    wire N__17123;
    wire N__17122;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17110;
    wire N__17105;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17095;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17076;
    wire N__17073;
    wire N__17066;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17040;
    wire N__17039;
    wire N__17038;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17022;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17010;
    wire N__17007;
    wire N__17006;
    wire N__17003;
    wire N__17002;
    wire N__16999;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16977;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16938;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16915;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16893;
    wire N__16890;
    wire N__16885;
    wire N__16884;
    wire N__16883;
    wire N__16882;
    wire N__16879;
    wire N__16878;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16864;
    wire N__16857;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16833;
    wire N__16832;
    wire N__16829;
    wire N__16828;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16821;
    wire N__16818;
    wire N__16817;
    wire N__16816;
    wire N__16813;
    wire N__16812;
    wire N__16811;
    wire N__16810;
    wire N__16807;
    wire N__16800;
    wire N__16795;
    wire N__16794;
    wire N__16791;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16768;
    wire N__16765;
    wire N__16760;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16728;
    wire N__16725;
    wire N__16724;
    wire N__16723;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16719;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16711;
    wire N__16710;
    wire N__16707;
    wire N__16706;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16695;
    wire N__16694;
    wire N__16689;
    wire N__16686;
    wire N__16685;
    wire N__16678;
    wire N__16675;
    wire N__16668;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16640;
    wire N__16633;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16607;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16568;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16512;
    wire N__16511;
    wire N__16510;
    wire N__16509;
    wire N__16506;
    wire N__16501;
    wire N__16492;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16487;
    wire N__16486;
    wire N__16485;
    wire N__16484;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16469;
    wire N__16464;
    wire N__16461;
    wire N__16456;
    wire N__16451;
    wire N__16448;
    wire N__16443;
    wire N__16438;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16409;
    wire N__16408;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16388;
    wire N__16387;
    wire N__16384;
    wire N__16383;
    wire N__16382;
    wire N__16379;
    wire N__16378;
    wire N__16375;
    wire N__16374;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16346;
    wire N__16343;
    wire N__16336;
    wire N__16329;
    wire N__16326;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16288;
    wire N__16285;
    wire N__16280;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16263;
    wire N__16262;
    wire N__16257;
    wire N__16256;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16252;
    wire N__16249;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16231;
    wire N__16230;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16218;
    wire N__16215;
    wire N__16214;
    wire N__16209;
    wire N__16206;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16108;
    wire N__16105;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16069;
    wire N__16064;
    wire N__16059;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15996;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15987;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15978;
    wire N__15977;
    wire N__15974;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15966;
    wire N__15961;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15893;
    wire N__15890;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15849;
    wire N__15848;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15836;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15795;
    wire N__15794;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15786;
    wire N__15785;
    wire N__15782;
    wire N__15773;
    wire N__15768;
    wire N__15765;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15738;
    wire N__15737;
    wire N__15736;
    wire N__15733;
    wire N__15728;
    wire N__15725;
    wire N__15720;
    wire N__15717;
    wire N__15716;
    wire N__15715;
    wire N__15714;
    wire N__15713;
    wire N__15712;
    wire N__15711;
    wire N__15708;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15688;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15676;
    wire N__15675;
    wire N__15674;
    wire N__15673;
    wire N__15672;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15654;
    wire N__15653;
    wire N__15652;
    wire N__15651;
    wire N__15644;
    wire N__15643;
    wire N__15642;
    wire N__15641;
    wire N__15640;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15620;
    wire N__15617;
    wire N__15612;
    wire N__15605;
    wire N__15598;
    wire N__15591;
    wire N__15582;
    wire N__15581;
    wire N__15580;
    wire N__15579;
    wire N__15578;
    wire N__15577;
    wire N__15574;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15543;
    wire N__15542;
    wire N__15541;
    wire N__15540;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15503;
    wire N__15496;
    wire N__15477;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15471;
    wire N__15470;
    wire N__15467;
    wire N__15460;
    wire N__15453;
    wire N__15452;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15434;
    wire N__15431;
    wire N__15430;
    wire N__15429;
    wire N__15428;
    wire N__15419;
    wire N__15416;
    wire N__15411;
    wire N__15408;
    wire N__15399;
    wire N__15398;
    wire N__15397;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15386;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15356;
    wire N__15353;
    wire N__15348;
    wire N__15339;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15332;
    wire N__15331;
    wire N__15330;
    wire N__15329;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15317;
    wire N__15314;
    wire N__15313;
    wire N__15312;
    wire N__15311;
    wire N__15310;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15292;
    wire N__15287;
    wire N__15284;
    wire N__15283;
    wire N__15282;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15274;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15262;
    wire N__15261;
    wire N__15260;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15245;
    wire N__15232;
    wire N__15229;
    wire N__15222;
    wire N__15215;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15193;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15188;
    wire N__15187;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15162;
    wire N__15159;
    wire N__15158;
    wire N__15157;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15149;
    wire N__15144;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15128;
    wire N__15125;
    wire N__15124;
    wire N__15119;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15082;
    wire N__15073;
    wire N__15054;
    wire N__15053;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15045;
    wire N__15044;
    wire N__15043;
    wire N__15040;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14990;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14983;
    wire N__14982;
    wire N__14981;
    wire N__14980;
    wire N__14979;
    wire N__14978;
    wire N__14977;
    wire N__14976;
    wire N__14975;
    wire N__14974;
    wire N__14967;
    wire N__14960;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14942;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14934;
    wire N__14927;
    wire N__14922;
    wire N__14919;
    wire N__14914;
    wire N__14903;
    wire N__14902;
    wire N__14901;
    wire N__14900;
    wire N__14897;
    wire N__14892;
    wire N__14887;
    wire N__14886;
    wire N__14883;
    wire N__14878;
    wire N__14873;
    wire N__14870;
    wire N__14863;
    wire N__14860;
    wire N__14855;
    wire N__14850;
    wire N__14847;
    wire N__14840;
    wire N__14837;
    wire N__14832;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14816;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14804;
    wire N__14803;
    wire N__14802;
    wire N__14799;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14786;
    wire N__14785;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14758;
    wire N__14753;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14732;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14684;
    wire N__14683;
    wire N__14682;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14670;
    wire N__14669;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14652;
    wire N__14651;
    wire N__14650;
    wire N__14649;
    wire N__14646;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14602;
    wire N__14589;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14529;
    wire N__14528;
    wire N__14527;
    wire N__14526;
    wire N__14525;
    wire N__14522;
    wire N__14521;
    wire N__14520;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14505;
    wire N__14504;
    wire N__14503;
    wire N__14498;
    wire N__14493;
    wire N__14488;
    wire N__14487;
    wire N__14486;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14470;
    wire N__14463;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14442;
    wire N__14437;
    wire N__14434;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14405;
    wire N__14400;
    wire N__14397;
    wire N__14396;
    wire N__14395;
    wire N__14394;
    wire N__14391;
    wire N__14390;
    wire N__14389;
    wire N__14388;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14384;
    wire N__14381;
    wire N__14376;
    wire N__14375;
    wire N__14374;
    wire N__14371;
    wire N__14362;
    wire N__14357;
    wire N__14354;
    wire N__14353;
    wire N__14352;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14340;
    wire N__14337;
    wire N__14332;
    wire N__14329;
    wire N__14328;
    wire N__14325;
    wire N__14320;
    wire N__14313;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14256;
    wire N__14255;
    wire N__14252;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14224;
    wire N__14217;
    wire N__14216;
    wire N__14213;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14197;
    wire N__14194;
    wire N__14181;
    wire N__14180;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14172;
    wire N__14167;
    wire N__14166;
    wire N__14163;
    wire N__14162;
    wire N__14161;
    wire N__14160;
    wire N__14155;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14125;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14103;
    wire N__14102;
    wire N__14101;
    wire N__14100;
    wire N__14099;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14085;
    wire N__14084;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14058;
    wire N__14057;
    wire N__14054;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14038;
    wire N__14033;
    wire N__14026;
    wire N__14021;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13985;
    wire N__13982;
    wire N__13981;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13966;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13919;
    wire N__13918;
    wire N__13917;
    wire N__13914;
    wire N__13913;
    wire N__13912;
    wire N__13909;
    wire N__13908;
    wire N__13905;
    wire N__13904;
    wire N__13901;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13851;
    wire N__13842;
    wire N__13833;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13812;
    wire N__13811;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13794;
    wire N__13787;
    wire N__13776;
    wire N__13773;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13767;
    wire N__13766;
    wire N__13763;
    wire N__13762;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13742;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13626;
    wire N__13623;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13586;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire N__13576;
    wire N__13569;
    wire N__13566;
    wire N__13565;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13548;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13539;
    wire N__13532;
    wire N__13531;
    wire N__13526;
    wire N__13523;
    wire N__13518;
    wire N__13517;
    wire N__13516;
    wire N__13511;
    wire N__13508;
    wire N__13507;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13499;
    wire N__13496;
    wire N__13489;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13458;
    wire N__13457;
    wire N__13456;
    wire N__13453;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13431;
    wire N__13428;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13410;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13389;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13293;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13261;
    wire N__13256;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13221;
    wire N__13218;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13183;
    wire N__13182;
    wire N__13179;
    wire N__13174;
    wire N__13171;
    wire N__13164;
    wire N__13163;
    wire N__13162;
    wire N__13159;
    wire N__13158;
    wire N__13155;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13131;
    wire N__13130;
    wire N__13127;
    wire N__13126;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13106;
    wire N__13103;
    wire N__13102;
    wire N__13099;
    wire N__13098;
    wire N__13095;
    wire N__13088;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13049;
    wire N__13048;
    wire N__13045;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13025;
    wire N__13018;
    wire N__13015;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12982;
    wire N__12973;
    wire N__12972;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12959;
    wire N__12954;
    wire N__12951;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12921;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12913;
    wire N__12912;
    wire N__12903;
    wire N__12902;
    wire N__12901;
    wire N__12898;
    wire N__12893;
    wire N__12890;
    wire N__12889;
    wire N__12888;
    wire N__12887;
    wire N__12884;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12872;
    wire N__12863;
    wire N__12858;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12804;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12777;
    wire N__12776;
    wire N__12773;
    wire N__12772;
    wire N__12771;
    wire N__12770;
    wire N__12763;
    wire N__12760;
    wire N__12759;
    wire N__12756;
    wire N__12755;
    wire N__12754;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12737;
    wire N__12736;
    wire N__12733;
    wire N__12732;
    wire N__12731;
    wire N__12728;
    wire N__12727;
    wire N__12722;
    wire N__12717;
    wire N__12710;
    wire N__12707;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12686;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12608;
    wire N__12607;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12595;
    wire N__12594;
    wire N__12591;
    wire N__12582;
    wire N__12577;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12513;
    wire N__12512;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12500;
    wire N__12495;
    wire N__12492;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12477;
    wire N__12476;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12448;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12434;
    wire N__12433;
    wire N__12432;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12426;
    wire N__12425;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12398;
    wire N__12391;
    wire N__12372;
    wire N__12369;
    wire N__12368;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12360;
    wire N__12359;
    wire N__12358;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12341;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12327;
    wire N__12326;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12303;
    wire N__12300;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12261;
    wire N__12258;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12246;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12217;
    wire N__12216;
    wire N__12215;
    wire N__12214;
    wire N__12213;
    wire N__12210;
    wire N__12209;
    wire N__12208;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12196;
    wire N__12193;
    wire N__12188;
    wire N__12181;
    wire N__12178;
    wire N__12173;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12147;
    wire N__12146;
    wire N__12143;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12120;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12064;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12052;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11947;
    wire N__11944;
    wire N__11943;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11919;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11861;
    wire N__11860;
    wire N__11857;
    wire N__11852;
    wire N__11847;
    wire N__11844;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11821;
    wire N__11818;
    wire N__11813;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11768;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11733;
    wire N__11732;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11715;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11692;
    wire N__11689;
    wire N__11684;
    wire N__11681;
    wire N__11674;
    wire N__11667;
    wire N__11666;
    wire N__11665;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11657;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11640;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11621;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11596;
    wire N__11591;
    wire N__11588;
    wire N__11583;
    wire N__11574;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11556;
    wire N__11551;
    wire N__11546;
    wire N__11541;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11525;
    wire N__11524;
    wire N__11521;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11503;
    wire N__11496;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11330;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11297;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11261;
    wire N__11252;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11226;
    wire N__11223;
    wire N__11222;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11168;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11156;
    wire N__11153;
    wire N__11152;
    wire N__11151;
    wire N__11142;
    wire N__11139;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11127;
    wire N__11122;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11103;
    wire N__11096;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11038;
    wire N__11033;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10910;
    wire N__10905;
    wire N__10902;
    wire N__10901;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10829;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10785;
    wire N__10776;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10759;
    wire N__10752;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10740;
    wire N__10739;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10722;
    wire N__10721;
    wire N__10718;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10702;
    wire N__10695;
    wire N__10694;
    wire N__10691;
    wire N__10686;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10659;
    wire N__10658;
    wire N__10657;
    wire N__10656;
    wire N__10653;
    wire N__10648;
    wire N__10645;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10631;
    wire N__10624;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10583;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10566;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10556;
    wire N__10553;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10509;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10430;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10413;
    wire N__10412;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10391;
    wire N__10390;
    wire N__10389;
    wire N__10388;
    wire N__10387;
    wire N__10384;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10362;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10339;
    wire N__10334;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10318;
    wire N__10311;
    wire N__10310;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10302;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10256;
    wire N__10255;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10172;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10160;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10135;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10109;
    wire N__10106;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10094;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10073;
    wire N__10070;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10059;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10041;
    wire N__10040;
    wire N__10039;
    wire N__10036;
    wire N__10031;
    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10021;
    wire N__10016;
    wire N__10011;
    wire N__10008;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9969;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9951;
    wire N__9948;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9888;
    wire N__9885;
    wire N__9884;
    wire N__9883;
    wire N__9880;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9868;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9827;
    wire N__9822;
    wire N__9815;
    wire N__9810;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9798;
    wire N__9797;
    wire N__9796;
    wire N__9795;
    wire N__9792;
    wire N__9785;
    wire N__9780;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9771;
    wire N__9768;
    wire N__9763;
    wire N__9760;
    wire N__9753;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9743;
    wire N__9738;
    wire N__9733;
    wire N__9726;
    wire N__9723;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9719;
    wire N__9716;
    wire N__9709;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9696;
    wire N__9691;
    wire N__9686;
    wire N__9679;
    wire N__9674;
    wire N__9663;
    wire N__9660;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9652;
    wire N__9647;
    wire N__9644;
    wire N__9643;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9599;
    wire N__9594;
    wire N__9591;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9579;
    wire N__9578;
    wire N__9573;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9507;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9405;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9386;
    wire N__9383;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9373;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9361;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9347;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9330;
    wire N__9329;
    wire N__9326;
    wire N__9325;
    wire N__9324;
    wire N__9321;
    wire N__9320;
    wire N__9317;
    wire N__9312;
    wire N__9309;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9297;
    wire N__9294;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9276;
    wire N__9265;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9259;
    wire N__9254;
    wire N__9245;
    wire N__9240;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9122;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9110;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9087;
    wire N__9084;
    wire N__9083;
    wire N__9078;
    wire N__9075;
    wire N__9074;
    wire N__9069;
    wire N__9066;
    wire N__9065;
    wire N__9064;
    wire N__9063;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9045;
    wire N__9042;
    wire N__9041;
    wire N__9038;
    wire N__9037;
    wire N__9034;
    wire N__9029;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9018;
    wire N__9011;
    wire N__9008;
    wire N__9003;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8982;
    wire N__8979;
    wire N__8978;
    wire N__8975;
    wire N__8974;
    wire N__8971;
    wire N__8966;
    wire N__8963;
    wire N__8958;
    wire N__8957;
    wire N__8952;
    wire N__8949;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8940;
    wire N__8937;
    wire N__8932;
    wire N__8929;
    wire N__8922;
    wire N__8921;
    wire N__8920;
    wire N__8919;
    wire N__8914;
    wire N__8913;
    wire N__8912;
    wire N__8907;
    wire N__8904;
    wire N__8899;
    wire N__8892;
    wire N__8889;
    wire N__8888;
    wire N__8887;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8874;
    wire N__8873;
    wire N__8872;
    wire N__8871;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8853;
    wire N__8850;
    wire N__8845;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8821;
    wire N__8818;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8787;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8775;
    wire N__8770;
    wire N__8767;
    wire N__8760;
    wire N__8757;
    wire N__8756;
    wire N__8755;
    wire N__8754;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8732;
    wire N__8727;
    wire N__8718;
    wire N__8715;
    wire N__8714;
    wire N__8711;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8697;
    wire N__8694;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8613;
    wire N__8612;
    wire N__8611;
    wire N__8606;
    wire N__8603;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8588;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8571;
    wire N__8568;
    wire N__8567;
    wire N__8566;
    wire N__8565;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8536;
    wire N__8533;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8513;
    wire N__8512;
    wire N__8511;
    wire N__8508;
    wire N__8503;
    wire N__8500;
    wire N__8495;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8351;
    wire N__8346;
    wire N__8343;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8331;
    wire N__8328;
    wire N__8327;
    wire N__8326;
    wire N__8325;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8311;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8292;
    wire N__8289;
    wire N__8288;
    wire N__8287;
    wire N__8284;
    wire N__8283;
    wire N__8282;
    wire N__8279;
    wire N__8274;
    wire N__8269;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8255;
    wire N__8254;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8228;
    wire N__8227;
    wire N__8224;
    wire N__8219;
    wire N__8216;
    wire N__8211;
    wire N__8208;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8174;
    wire N__8173;
    wire N__8170;
    wire N__8165;
    wire N__8162;
    wire N__8157;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8151;
    wire N__8150;
    wire N__8141;
    wire N__8138;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8123;
    wire N__8120;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8109;
    wire N__8100;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8092;
    wire N__8081;
    wire N__8078;
    wire N__8073;
    wire N__8070;
    wire N__8069;
    wire N__8068;
    wire N__8067;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8051;
    wire N__8046;
    wire N__8043;
    wire N__8042;
    wire N__8041;
    wire N__8040;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8012;
    wire N__8011;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8005;
    wire N__7992;
    wire N__7989;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7940;
    wire N__7939;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7923;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7896;
    wire N__7895;
    wire N__7894;
    wire N__7891;
    wire N__7890;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7886;
    wire N__7881;
    wire N__7876;
    wire N__7871;
    wire N__7868;
    wire N__7859;
    wire N__7854;
    wire N__7845;
    wire N__7844;
    wire N__7841;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7829;
    wire N__7824;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7812;
    wire N__7811;
    wire N__7810;
    wire N__7807;
    wire N__7802;
    wire N__7797;
    wire N__7794;
    wire N__7793;
    wire N__7790;
    wire N__7789;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7777;
    wire N__7774;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7742;
    wire N__7741;
    wire N__7738;
    wire N__7737;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7716;
    wire N__7715;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7705;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7689;
    wire N__7686;
    wire N__7685;
    wire N__7684;
    wire N__7683;
    wire N__7682;
    wire N__7679;
    wire N__7674;
    wire N__7669;
    wire N__7664;
    wire N__7659;
    wire N__7656;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7634;
    wire N__7631;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7595;
    wire N__7592;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7572;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7564;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7552;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7461;
    wire N__7458;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7344;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7326;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7304;
    wire N__7301;
    wire N__7300;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7288;
    wire N__7281;
    wire N__7280;
    wire N__7279;
    wire N__7276;
    wire N__7271;
    wire N__7268;
    wire N__7263;
    wire N__7262;
    wire N__7261;
    wire N__7260;
    wire N__7257;
    wire N__7256;
    wire N__7247;
    wire N__7244;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7209;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7203;
    wire N__7196;
    wire N__7193;
    wire N__7188;
    wire N__7187;
    wire N__7186;
    wire N__7183;
    wire N__7178;
    wire N__7175;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu2.r_data_wire_4 ;
    wire \INVuu2.r_data_reg_4C_net ;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \uu0.un88_ci_3_cascade_ ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.un4_l_count_13_cascade_ ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.un11_l_count_i ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.un4_l_count_16 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un66_ci ;
    wire \uu0.un88_ci_3 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.r_data_wire_0 ;
    wire vbuf_tx_data_0;
    wire \uu2.r_data_wire_1 ;
    wire vbuf_tx_data_1;
    wire \uu2.r_data_wire_2 ;
    wire vbuf_tx_data_2;
    wire \uu2.r_data_wire_3 ;
    wire vbuf_tx_data_3;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.un404_ci_cascade_ ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.un165_ci_0 ;
    wire \uu0.sec_clkDZ0 ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.un404_ci ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \INVuu2.bitmap_111C_net ;
    wire \uu0.un55_ci ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.un110_ci ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \buart.Z_tx.un1_bitcount_c3_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \Lab_UT.alarmchar10_i_2 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_2 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_6 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_7 ;
    wire \uu2.N_102_cascade_ ;
    wire \uu2.N_61_i ;
    wire \INVuu2.w_addr_user_8C_net ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_4 ;
    wire \uu2.w_addr_user_3_i_a2_3_6 ;
    wire \uu2.mem0.g1_3_0_cascade_ ;
    wire \uu2.mem0.N_63_0_i ;
    wire \uu2.mem0.G_17_0_0_0 ;
    wire N_72_mux;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_3 ;
    wire \uu2.w_addr_user_3_i_a2_2_6 ;
    wire \uu2.un28_w_addr_user_i_0_cascade_ ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.N_105 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \INVuu2.w_addr_user_1C_net ;
    wire \uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_ ;
    wire \Lab_UT.alarmchar_2_1_1 ;
    wire \resetGen.reset_count_2_0_4_cascade_ ;
    wire \Lab_UT.alarmchar10 ;
    wire \Lab_UT.alarmcharZ0Z_4 ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.un241_ci ;
    wire \resetGen.un241_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire vbuf_tx_data_rdy;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.un143_ci_0 ;
    wire \uu2.un1_l_count_1_2_0_cascade_ ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu2.un1_l_count_2_2_cascade_ ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire bfn_4_13_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.ser_clk ;
    wire \uu2.N_155 ;
    wire \uu2.N_106 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.N_102 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.N_97 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \INVuu2.w_addr_user_nesr_0C_net ;
    wire \uu2.un28_w_addr_user_i_0_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_12 ;
    wire \uu2.N_41_0_cascade_ ;
    wire \uu2.N_132_mux ;
    wire \uu2.N_132_mux_cascade_ ;
    wire \uu2.mem0.N_94_i ;
    wire \uu2.N_15_i ;
    wire \uu2.un21_w_addr_displaying_i_cascade_ ;
    wire \INVuu2.w_addr_displaying_0C_net ;
    wire \Lab_UT.alarmcharZ0Z_5 ;
    wire \uu2.mem0.N_13_1_0_0 ;
    wire \uu2.mem0.i14_mux_0_0_0_cascade_ ;
    wire \uu2.mem0.N_8_0_0_1 ;
    wire \Lab_UT.alarmcharZ0Z_6 ;
    wire \Lab_UT.bcd2segment1.m68_bmZ0 ;
    wire \uu2.un28_w_addr_user_i_0_a2Z0Z_4 ;
    wire L3_tx_data_3;
    wire L3_tx_data_4;
    wire L3_tx_data_0;
    wire \uu2.w_data_i_o2_4Z0Z_0_cascade_ ;
    wire N_96_cascade_;
    wire \Lab_UT.bcd2segment1.m59_bmZ0 ;
    wire \Lab_UT.bcd2segment1.m52_amZ0 ;
    wire \Lab_UT.alarmcharZ0Z_0 ;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z_0 ;
    wire \Lab_UT.dictrl.next_alarmstate_1 ;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_ ;
    wire \Lab_UT.bcd2segment1.m59_amZ0 ;
    wire \Lab_UT.dictrl.un1_next_alarmstate21_0 ;
    wire \Lab_UT.cnt_0 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu0.un4_l_count_0 ;
    wire o_One_Sec_Pulse;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu2.un284_ci ;
    wire \uu2.l_countZ0Z_2 ;
    wire uart_RXD;
    wire \uu2.un350_ci ;
    wire \uu2.l_countZ0Z_8 ;
    wire \Lab_UT.dictrl.next_alarmstate_0_0 ;
    wire \Lab_UT.dictrl.G_74 ;
    wire \Lab_UT.bcd2segment1.N_187_cascade_ ;
    wire \Lab_UT.bcd2segment1.N_189_cascade_ ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.mem0.N_107_0_cascade_ ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_1 ;
    wire L3_tx_data_6;
    wire \uu2.mem0.N_130_mux_cascade_ ;
    wire \uu2.mem0.N_54_0_i ;
    wire \uu2.mem0.N_17_0_cascade_ ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_5 ;
    wire \uu2.mem0.N_107_0_0 ;
    wire \uu2.mem0.N_74_0_0_1 ;
    wire \uu2.mem0.g0_7_0_0_2_cascade_ ;
    wire \uu2.mem0.N_3_0_cascade_ ;
    wire \uu2.mem0.N_98_0_0_0 ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \uu2.N_1585_0_0 ;
    wire \Lab_UT.bcd2segment1.i6_mux_cascade_ ;
    wire \Lab_UT.bcd2segment1.m68_amZ0 ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire rst;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_0 ;
    wire clk;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_ ;
    wire \uu2.mem0.g1_2_0 ;
    wire \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0 ;
    wire \uu2.mem0.g0_7_0_0_1 ;
    wire \INVuu2.w_addr_displaying_nesr_3C_net ;
    wire \Lab_UT.alarmchar9_cascade_ ;
    wire \Lab_UT.alarmcharZ0Z_2 ;
    wire \Lab_UT.bcd2segment1.N_160 ;
    wire \Lab_UT.bcd2segment1.i5_mux_cascade_ ;
    wire \Lab_UT.cnt_2 ;
    wire \Lab_UT.bcd2segment1.m42_amZ0_cascade_ ;
    wire \Lab_UT.bcd2segment1.m52_bmZ0 ;
    wire \Lab_UT.bcd2segment1.N_42_i ;
    wire \Lab_UT.dictrl.alarmstateZ0Z_0 ;
    wire \Lab_UT.dictrl.idle_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstate_1_0 ;
    wire \Lab_UT.bcd2segment1.N_222_cascade_ ;
    wire \Lab_UT.dictrl.alarmstateZ0Z_1 ;
    wire \Lab_UT.dictrl.alarmstate_i_3_0 ;
    wire \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \Lab_UT.q_5_1_cascade_ ;
    wire \buart.Z_rx.ser_clk_2_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z4 ;
    wire \Lab_UT.dictrl.next_alarmstate4Z0Z_0 ;
    wire \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0 ;
    wire \Lab_UT.bcd2segment1.N_194_cascade_ ;
    wire \uu2.mem0.N_92_0_cascade_ ;
    wire \uu2.mem0.m73_ns_1_0 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_1_4 ;
    wire \INVuu2.bitmap_90C_net ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.mem0.N_92_0_0_cascade_ ;
    wire \uu2.mem0.m73_ns_1_0_0_1 ;
    wire \uu2.mem0.N_74_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_34 ;
    wire L3_tx_data_2;
    wire \uu2.mem0.N_93_i ;
    wire \uu2.mem0.N_57_0_0 ;
    wire \uu2.mem0.N_67_0 ;
    wire \uu2.mem0.g0_1_cascade_ ;
    wire \uu2.mem0.g0_2 ;
    wire \uu2.mem0.i14_mux ;
    wire \uu2.mem0.N_126_0 ;
    wire \uu2.mem0.g0_1_3_cascade_ ;
    wire \uu2.mem0.G_13_0_a2_0_1 ;
    wire \uu2.mem0.N_22_cascade_ ;
    wire \uu2.mem0.N_66_0_i ;
    wire \uu2.mem0.g0_i_m2_1 ;
    wire \uu2.mem0.g2_0_0_0 ;
    wire \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1 ;
    wire \uu2.N_67_1_0 ;
    wire \uu2.N_67_1_0_cascade_ ;
    wire \uu2.mem0.N_55_0_0_0 ;
    wire \uu2.mem0.g2_1 ;
    wire \INVuu2.w_addr_displaying_1C_net ;
    wire \Lab_UT.bcd2segment1.N_250_cascade_ ;
    wire \Lab_UT.bcd2segment1.i2_mux_cascade_ ;
    wire \INVuu2.bitmap_296C_net ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.m95_i_m2_i_m2_1_cascade_ ;
    wire \uu2.N_16_cascade_ ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_3_rep1_nesrC_net ;
    wire \Lab_UT.N_27_i ;
    wire \resetGen.escKeyZ0Z_4 ;
    wire \resetGen.escKeyZ0 ;
    wire \Lab_UT.didp.did_alarmMatch_1_cascade_ ;
    wire \Lab_UT.zero ;
    wire \Lab_UT.alarmMatch ;
    wire \Lab_UT.didp.countrce3.did_alarmMatch_0 ;
    wire \Lab_UT.q_5_3 ;
    wire \Lab_UT.q_5_0_cascade_ ;
    wire \Lab_UT.q_5_2 ;
    wire \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.next_state_out_1 ;
    wire \Lab_UT.dictrl.N_97_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_7_12_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa_1 ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_ ;
    wire \resetGen.escKeyZ0Z_5 ;
    wire \Lab_UT.dictrl.next_state_set_0_1 ;
    wire bu_rx_data_6;
    wire bu_rx_data_7;
    wire bu_rx_data_4;
    wire \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0 ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5 ;
    wire \Lab_UT.dictrl.un1_state_16_cascade_ ;
    wire bu_rx_data_5;
    wire bu_rx_data_1;
    wire bu_rx_data_0;
    wire \Lab_UT.bcd2segment1.N_127_mux_cascade_ ;
    wire \Lab_UT.bcd2segment1.N_235_cascade_ ;
    wire \Lab_UT.bcd2segment1.N_237_cascade_ ;
    wire \INVuu2.bitmap_162C_net ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.N_101_0 ;
    wire \Lab_UT.bcd2segment1.N_242_cascade_ ;
    wire \Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_ ;
    wire \uu2.N_1580_0_cascade_ ;
    wire \uu2.N_77_0 ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.N_1581_0 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \INVuu2.bitmap_75C_net ;
    wire L3_tx_data_5;
    wire \uu2.mem0.N_134_mux_cascade_ ;
    wire \uu2.w_data_i_0_tzZ0Z_0 ;
    wire \uu2.mem0.N_60_0_i ;
    wire \uu2.mem0.N_55_0 ;
    wire \uu2.N_126_cascade_ ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_67 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_66 ;
    wire \uu2.N_126 ;
    wire \uu2.mem0.g0_7_0_0 ;
    wire \uu2.mem0.N_57_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_u_i_5_1 ;
    wire \uu2.mem0.g0_7_0_3 ;
    wire \uu2.N_16 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_57 ;
    wire \uu2.mem0.N_13_0 ;
    wire \uu2.N_8 ;
    wire \uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8 ;
    wire \uu2.w_addr_displaying_fastZ0Z_4 ;
    wire \INVuu2.w_addr_displaying_4_rep1C_net ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.N_9_i ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \uu2.mem0.N_9_cascade_ ;
    wire \uu2.mem0.N_15 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.mem0.N_7 ;
    wire \uu2.mem0.m317_0_a6_0_cascade_ ;
    wire \uu2.mem0.N_6_0 ;
    wire \uu2.mem0.m317_0_0 ;
    wire \uu2.mem0.N_11_0_0_cascade_ ;
    wire \uu2.mem0.N_6_0_0_0 ;
    wire \uu2.w_addr_displaying_4_repZ0Z1 ;
    wire \uu2.mem0.N_5_0 ;
    wire \uu2.mem0.N_14 ;
    wire \uu2.mem0.g1_2_2_2_1 ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \Lab_UT.bcd2segment1.N_239 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.N_115 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \INVuu2.bitmap_34C_net ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_ ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_0 ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_ ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \INVuu2.bitmap_180C_net ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_ ;
    wire \Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.N_9_0 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.bcd2segment1.N_181 ;
    wire \Lab_UT.bcd2segment1.N_229 ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.bcd2segment1.N_233 ;
    wire \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1 ;
    wire \Lab_UT.dictrl.dicRun_2_reti ;
    wire \Lab_UT.dictrl.next_state_out_0 ;
    wire \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ;
    wire \Lab_UT.dictrl.next_state_set ;
    wire \buart.Z_rx.bitcount_lm_3_cascade_ ;
    wire \Lab_UT.m72_0 ;
    wire \Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1 ;
    wire \Lab_UT.un1_state_13 ;
    wire \Lab_UT.un1_state_13_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \Lab_UT.dictrl.un1_state_11 ;
    wire \Lab_UT.dictrl.un1_state_11_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1 ;
    wire \Lab_UT.bcd2segment1.N_264 ;
    wire \Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.next_state16Z0Z_5 ;
    wire \Lab_UT.m68_0_ns_cascade_ ;
    wire \Lab_UT.dictrl.next_state16Z0Z_4 ;
    wire \Lab_UT.state_3 ;
    wire \Lab_UT.state_1 ;
    wire \Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_ ;
    wire \Lab_UT.state_2 ;
    wire \Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_1 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.m76_am_1 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \Lab_UT.bcd2segment1.N_244 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \Lab_UT.bcd2segment1.N_246_cascade_ ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.di_Mones_3 ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.bcd2segment1.N_248_cascade_ ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.m76_bm_1_0 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \INVuu2.bitmap_168C_net ;
    wire \uu2.mem0.g1_2_2 ;
    wire \uu2.mem0.g2_0_0_0_0 ;
    wire \uu2.mem0.g2_2 ;
    wire \uu2.w_addr_displaying_2_repZ0Z1 ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_u_i_4_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_69 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \INVuu2.w_addr_displaying_ness_6C_net ;
    wire \uu2.un21_w_addr_displaying_i_0 ;
    wire \uu2.mem0.G_13_0_a2_1_cascade_ ;
    wire \uu2.mem0.G_13_0_a3_1_2 ;
    wire L3_tx_data_rdy;
    wire L3_tx_data_1;
    wire \uu2.mem0.G_13_0_a2_2_cascade_ ;
    wire N_96;
    wire \uu2.mem0.G_13_0_0 ;
    wire \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0 ;
    wire \uu2.N_12_i_cascade_ ;
    wire \uu2.N_67 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.un21_w_addr_displaying_i ;
    wire \uu2.N_12_i ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \INVuu2.w_addr_displaying_7_rep1C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.N_272_cascade_ ;
    wire \uu2.mem0.m317_0_a6_1_0 ;
    wire \uu2.mem0.N_13 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \Lab_UT.Run ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \INVuu2.bitmap_58C_net ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.w_addr_displaying_8_repZ0Z1 ;
    wire \uu2.N_272 ;
    wire \uu2.w_addr_displaying_3_repZ0Z2 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_ ;
    wire \uu2.mem0.N_294 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.mem0.N_271 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_80 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.w_addr_displaying_7_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \uu2.mem0.N_98_0 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.bcd2segment1.N_166 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.didp.countrce3.q_RNO_0Z0Z_3 ;
    wire bfn_9_10_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcount_lm_4 ;
    wire \Lab_UT.alarmcharZ0Z_1 ;
    wire \Lab_UT.cnt_3 ;
    wire \Lab_UT.cnt_1 ;
    wire \Lab_UT.bcd2segment1.m42_bmZ0 ;
    wire CONSTANT_ONE_NET;
    wire \buart.Z_rx.bitcount_lm_0 ;
    wire \buart.Z_rx.un1_sample_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_out_3 ;
    wire \Lab_UT.m68_0_ns ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_lm_1 ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_lm_2 ;
    wire \Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ;
    wire \Lab_UT.dictrl.next_state_set_1 ;
    wire \Lab_UT.dictrl.un1_state_21_reti_i ;
    wire \Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2 ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \buart.Z_rx.valid_0_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire bu_rx_data_rdy_cascade_;
    wire \buart.Z_rx.N_27_0_i ;
    wire \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1 ;
    wire \Lab_UT.dictrl.next_state_out_2 ;
    wire \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \buart.Z_rx.idle_0 ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.ser_clk_2 ;
    wire \buart.Z_rx.ser_clk_3 ;
    wire \buart.Z_rx.idle_cascade_ ;
    wire bu_rx_data_rdy;
    wire \buart.Z_rx.bitcountlde_0 ;
    wire \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ;
    wire \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ;
    wire \Lab_UT.dictrl.next_state_set_2 ;
    wire \Lab_UT.state_i_3_3 ;
    wire \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ;
    wire \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1 ;
    wire \Lab_UT.dictrl.state_retZ0Z_4 ;
    wire \Lab_UT.dictrl.next_state_set_0 ;
    wire \Lab_UT.state_i_3_1 ;
    wire bu_rx_data_3;
    wire bu_rx_data_2;
    wire \buart.Z_rx.sample ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_0 ;
    wire \Lab_UT.bcd2segment1.N_192 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_5 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_3 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_4 ;
    wire \Lab_UT.three_2_cascade_ ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.didp.countrce2.un15_ce_2 ;
    wire \Lab_UT.didp.countrce2.un15_ce_2_cascade_ ;
    wire \Lab_UT.di_Stens_0 ;
    wire \Lab_UT.didp.countrce2.un20_qPone_cascade_ ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.three_2_0 ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.dictrl.dicRun_2 ;
    wire \Lab_UT.state_i_3_2 ;
    wire \Lab_UT.state_0 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.nine ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.q_RNI84NN1_2 ;
    wire rst_g;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire _gnd_net_;
    wire clk_g;
    wire oneSecStrb_i;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__7023),
            .RESETB(N__16614),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__7230,N__7599,N__7572,N__7746,N__7689,N__7638,N__15894,N__15764,N__15848}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__8394,N__8403,N__10212,N__8478,N__8433,N__8412,N__10128,N__10548,N__12111}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__10086,dangling_wire_31,N__11808,dangling_wire_32,N__9192,dangling_wire_33,N__8460,dangling_wire_34,N__11028,dangling_wire_35,N__10968,dangling_wire_36,N__9171}),
            .RCLKE(),
            .RCLK(N__18496),
            .RE(N__16607),
            .WCLKE(N__10508),
            .WCLK(N__18495),
            .WE(N__10509));
    IO_PAD led_obuft_3_iopad (
            .OE(N__19573),
            .DIN(N__19572),
            .DOUT(N__19571),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__19573),
            .PADOUT(N__19572),
            .PADIN(N__19571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__19564),
            .DIN(N__19563),
            .DOUT(N__19562),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__19564),
            .PADOUT(N__19563),
            .PADIN(N__19562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__19555),
            .DIN(N__19554),
            .DOUT(N__19553),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__19555),
            .PADOUT(N__19554),
            .PADIN(N__19553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__19546),
            .DIN(N__19545),
            .DOUT(N__19544),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__19546),
            .PADOUT(N__19545),
            .PADIN(N__19544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__19537),
            .DIN(N__19536),
            .DOUT(N__19535),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__19537),
            .PADOUT(N__19536),
            .PADIN(N__19535),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__18469),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__19528),
            .DIN(N__19527),
            .DOUT(N__19526),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__19528),
            .PADOUT(N__19527),
            .PADIN(N__19526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__19519),
            .DIN(N__19518),
            .DOUT(N__19517),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__19519),
            .PADOUT(N__19518),
            .PADIN(N__19517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__19510),
            .DIN(N__19509),
            .DOUT(N__19508),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__19510),
            .PADOUT(N__19509),
            .PADIN(N__19508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__19501),
            .DIN(N__19500),
            .DOUT(N__19499),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__19501),
            .PADOUT(N__19500),
            .PADIN(N__19499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__19492),
            .DIN(N__19491),
            .DOUT(N__19490),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__19492),
            .PADOUT(N__19491),
            .PADIN(N__19490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7038),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__4752 (
            .O(N__19473),
            .I(N__19469));
    InMux I__4751 (
            .O(N__19472),
            .I(N__19458));
    InMux I__4750 (
            .O(N__19469),
            .I(N__19458));
    InMux I__4749 (
            .O(N__19468),
            .I(N__19458));
    InMux I__4748 (
            .O(N__19467),
            .I(N__19458));
    LocalMux I__4747 (
            .O(N__19458),
            .I(N__19455));
    Odrv4 I__4746 (
            .O(N__19455),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__4745 (
            .O(N__19452),
            .I(N__19446));
    InMux I__4744 (
            .O(N__19451),
            .I(N__19446));
    LocalMux I__4743 (
            .O(N__19446),
            .I(\Lab_UT.three_2_0 ));
    InMux I__4742 (
            .O(N__19443),
            .I(N__19440));
    LocalMux I__4741 (
            .O(N__19440),
            .I(N__19437));
    Span4Mux_h I__4740 (
            .O(N__19437),
            .I(N__19425));
    InMux I__4739 (
            .O(N__19436),
            .I(N__19417));
    InMux I__4738 (
            .O(N__19435),
            .I(N__19417));
    InMux I__4737 (
            .O(N__19434),
            .I(N__19414));
    InMux I__4736 (
            .O(N__19433),
            .I(N__19407));
    InMux I__4735 (
            .O(N__19432),
            .I(N__19407));
    InMux I__4734 (
            .O(N__19431),
            .I(N__19407));
    InMux I__4733 (
            .O(N__19430),
            .I(N__19400));
    InMux I__4732 (
            .O(N__19429),
            .I(N__19400));
    InMux I__4731 (
            .O(N__19428),
            .I(N__19400));
    Span4Mux_h I__4730 (
            .O(N__19425),
            .I(N__19397));
    InMux I__4729 (
            .O(N__19424),
            .I(N__19390));
    InMux I__4728 (
            .O(N__19423),
            .I(N__19390));
    InMux I__4727 (
            .O(N__19422),
            .I(N__19390));
    LocalMux I__4726 (
            .O(N__19417),
            .I(N__19387));
    LocalMux I__4725 (
            .O(N__19414),
            .I(N__19382));
    LocalMux I__4724 (
            .O(N__19407),
            .I(N__19382));
    LocalMux I__4723 (
            .O(N__19400),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv4 I__4722 (
            .O(N__19397),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__4721 (
            .O(N__19390),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv12 I__4720 (
            .O(N__19387),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv12 I__4719 (
            .O(N__19382),
            .I(\Lab_UT.di_Stens_2 ));
    CascadeMux I__4718 (
            .O(N__19371),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    InMux I__4717 (
            .O(N__19368),
            .I(N__19364));
    InMux I__4716 (
            .O(N__19367),
            .I(N__19359));
    LocalMux I__4715 (
            .O(N__19364),
            .I(N__19356));
    InMux I__4714 (
            .O(N__19363),
            .I(N__19351));
    InMux I__4713 (
            .O(N__19362),
            .I(N__19351));
    LocalMux I__4712 (
            .O(N__19359),
            .I(N__19345));
    Span4Mux_v I__4711 (
            .O(N__19356),
            .I(N__19340));
    LocalMux I__4710 (
            .O(N__19351),
            .I(N__19340));
    InMux I__4709 (
            .O(N__19350),
            .I(N__19335));
    InMux I__4708 (
            .O(N__19349),
            .I(N__19330));
    InMux I__4707 (
            .O(N__19348),
            .I(N__19330));
    Span4Mux_v I__4706 (
            .O(N__19345),
            .I(N__19324));
    Span4Mux_h I__4705 (
            .O(N__19340),
            .I(N__19324));
    InMux I__4704 (
            .O(N__19339),
            .I(N__19319));
    InMux I__4703 (
            .O(N__19338),
            .I(N__19319));
    LocalMux I__4702 (
            .O(N__19335),
            .I(N__19314));
    LocalMux I__4701 (
            .O(N__19330),
            .I(N__19314));
    InMux I__4700 (
            .O(N__19329),
            .I(N__19309));
    Span4Mux_v I__4699 (
            .O(N__19324),
            .I(N__19306));
    LocalMux I__4698 (
            .O(N__19319),
            .I(N__19301));
    Span12Mux_s10_h I__4697 (
            .O(N__19314),
            .I(N__19301));
    InMux I__4696 (
            .O(N__19313),
            .I(N__19296));
    InMux I__4695 (
            .O(N__19312),
            .I(N__19296));
    LocalMux I__4694 (
            .O(N__19309),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__4693 (
            .O(N__19306),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv12 I__4692 (
            .O(N__19301),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__4691 (
            .O(N__19296),
            .I(\Lab_UT.di_Sones_2 ));
    InMux I__4690 (
            .O(N__19287),
            .I(N__19278));
    InMux I__4689 (
            .O(N__19286),
            .I(N__19275));
    InMux I__4688 (
            .O(N__19285),
            .I(N__19270));
    InMux I__4687 (
            .O(N__19284),
            .I(N__19270));
    InMux I__4686 (
            .O(N__19283),
            .I(N__19265));
    InMux I__4685 (
            .O(N__19282),
            .I(N__19265));
    InMux I__4684 (
            .O(N__19281),
            .I(N__19261));
    LocalMux I__4683 (
            .O(N__19278),
            .I(N__19257));
    LocalMux I__4682 (
            .O(N__19275),
            .I(N__19253));
    LocalMux I__4681 (
            .O(N__19270),
            .I(N__19250));
    LocalMux I__4680 (
            .O(N__19265),
            .I(N__19247));
    CascadeMux I__4679 (
            .O(N__19264),
            .I(N__19244));
    LocalMux I__4678 (
            .O(N__19261),
            .I(N__19240));
    InMux I__4677 (
            .O(N__19260),
            .I(N__19237));
    Span4Mux_v I__4676 (
            .O(N__19257),
            .I(N__19234));
    InMux I__4675 (
            .O(N__19256),
            .I(N__19231));
    Span4Mux_h I__4674 (
            .O(N__19253),
            .I(N__19228));
    Span4Mux_h I__4673 (
            .O(N__19250),
            .I(N__19221));
    Span4Mux_s3_v I__4672 (
            .O(N__19247),
            .I(N__19221));
    InMux I__4671 (
            .O(N__19244),
            .I(N__19218));
    InMux I__4670 (
            .O(N__19243),
            .I(N__19215));
    Span4Mux_h I__4669 (
            .O(N__19240),
            .I(N__19212));
    LocalMux I__4668 (
            .O(N__19237),
            .I(N__19203));
    Span4Mux_h I__4667 (
            .O(N__19234),
            .I(N__19203));
    LocalMux I__4666 (
            .O(N__19231),
            .I(N__19203));
    Span4Mux_v I__4665 (
            .O(N__19228),
            .I(N__19203));
    InMux I__4664 (
            .O(N__19227),
            .I(N__19198));
    InMux I__4663 (
            .O(N__19226),
            .I(N__19198));
    Span4Mux_h I__4662 (
            .O(N__19221),
            .I(N__19195));
    LocalMux I__4661 (
            .O(N__19218),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__4660 (
            .O(N__19215),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__4659 (
            .O(N__19212),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__4658 (
            .O(N__19203),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__4657 (
            .O(N__19198),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__4656 (
            .O(N__19195),
            .I(\Lab_UT.di_Sones_1 ));
    CascadeMux I__4655 (
            .O(N__19182),
            .I(N__19174));
    CascadeMux I__4654 (
            .O(N__19181),
            .I(N__19170));
    CascadeMux I__4653 (
            .O(N__19180),
            .I(N__19167));
    CascadeMux I__4652 (
            .O(N__19179),
            .I(N__19164));
    CascadeMux I__4651 (
            .O(N__19178),
            .I(N__19161));
    CascadeMux I__4650 (
            .O(N__19177),
            .I(N__19158));
    InMux I__4649 (
            .O(N__19174),
            .I(N__19155));
    InMux I__4648 (
            .O(N__19173),
            .I(N__19152));
    InMux I__4647 (
            .O(N__19170),
            .I(N__19147));
    InMux I__4646 (
            .O(N__19167),
            .I(N__19147));
    InMux I__4645 (
            .O(N__19164),
            .I(N__19142));
    InMux I__4644 (
            .O(N__19161),
            .I(N__19142));
    InMux I__4643 (
            .O(N__19158),
            .I(N__19137));
    LocalMux I__4642 (
            .O(N__19155),
            .I(N__19133));
    LocalMux I__4641 (
            .O(N__19152),
            .I(N__19130));
    LocalMux I__4640 (
            .O(N__19147),
            .I(N__19125));
    LocalMux I__4639 (
            .O(N__19142),
            .I(N__19125));
    CascadeMux I__4638 (
            .O(N__19141),
            .I(N__19122));
    CascadeMux I__4637 (
            .O(N__19140),
            .I(N__19119));
    LocalMux I__4636 (
            .O(N__19137),
            .I(N__19116));
    CascadeMux I__4635 (
            .O(N__19136),
            .I(N__19112));
    Span4Mux_h I__4634 (
            .O(N__19133),
            .I(N__19109));
    Span4Mux_v I__4633 (
            .O(N__19130),
            .I(N__19104));
    Span4Mux_v I__4632 (
            .O(N__19125),
            .I(N__19104));
    InMux I__4631 (
            .O(N__19122),
            .I(N__19099));
    InMux I__4630 (
            .O(N__19119),
            .I(N__19099));
    Span4Mux_h I__4629 (
            .O(N__19116),
            .I(N__19096));
    InMux I__4628 (
            .O(N__19115),
            .I(N__19091));
    InMux I__4627 (
            .O(N__19112),
            .I(N__19091));
    Span4Mux_v I__4626 (
            .O(N__19109),
            .I(N__19088));
    Span4Mux_h I__4625 (
            .O(N__19104),
            .I(N__19083));
    LocalMux I__4624 (
            .O(N__19099),
            .I(N__19083));
    Odrv4 I__4623 (
            .O(N__19096),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__4622 (
            .O(N__19091),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv4 I__4621 (
            .O(N__19088),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv4 I__4620 (
            .O(N__19083),
            .I(\Lab_UT.di_Sones_3 ));
    InMux I__4619 (
            .O(N__19074),
            .I(N__19065));
    InMux I__4618 (
            .O(N__19073),
            .I(N__19060));
    InMux I__4617 (
            .O(N__19072),
            .I(N__19060));
    InMux I__4616 (
            .O(N__19071),
            .I(N__19055));
    InMux I__4615 (
            .O(N__19070),
            .I(N__19055));
    InMux I__4614 (
            .O(N__19069),
            .I(N__19048));
    InMux I__4613 (
            .O(N__19068),
            .I(N__19048));
    LocalMux I__4612 (
            .O(N__19065),
            .I(N__19045));
    LocalMux I__4611 (
            .O(N__19060),
            .I(N__19040));
    LocalMux I__4610 (
            .O(N__19055),
            .I(N__19040));
    InMux I__4609 (
            .O(N__19054),
            .I(N__19032));
    InMux I__4608 (
            .O(N__19053),
            .I(N__19032));
    LocalMux I__4607 (
            .O(N__19048),
            .I(N__19029));
    Span4Mux_s3_v I__4606 (
            .O(N__19045),
            .I(N__19026));
    Span4Mux_s3_v I__4605 (
            .O(N__19040),
            .I(N__19021));
    InMux I__4604 (
            .O(N__19039),
            .I(N__19014));
    InMux I__4603 (
            .O(N__19038),
            .I(N__19014));
    InMux I__4602 (
            .O(N__19037),
            .I(N__19014));
    LocalMux I__4601 (
            .O(N__19032),
            .I(N__19011));
    Span4Mux_v I__4600 (
            .O(N__19029),
            .I(N__19006));
    Span4Mux_v I__4599 (
            .O(N__19026),
            .I(N__19006));
    InMux I__4598 (
            .O(N__19025),
            .I(N__19001));
    InMux I__4597 (
            .O(N__19024),
            .I(N__19001));
    Span4Mux_h I__4596 (
            .O(N__19021),
            .I(N__18998));
    LocalMux I__4595 (
            .O(N__19014),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__4594 (
            .O(N__19011),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__4593 (
            .O(N__19006),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__4592 (
            .O(N__19001),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__4591 (
            .O(N__18998),
            .I(\Lab_UT.di_Sones_0 ));
    InMux I__4590 (
            .O(N__18987),
            .I(N__18984));
    LocalMux I__4589 (
            .O(N__18984),
            .I(N__18980));
    InMux I__4588 (
            .O(N__18983),
            .I(N__18977));
    Span12Mux_s1_h I__4587 (
            .O(N__18980),
            .I(N__18972));
    LocalMux I__4586 (
            .O(N__18977),
            .I(N__18972));
    Odrv12 I__4585 (
            .O(N__18972),
            .I(\Lab_UT.dictrl.dicRun_2 ));
    InMux I__4584 (
            .O(N__18969),
            .I(N__18964));
    InMux I__4583 (
            .O(N__18968),
            .I(N__18961));
    CascadeMux I__4582 (
            .O(N__18967),
            .I(N__18956));
    LocalMux I__4581 (
            .O(N__18964),
            .I(N__18949));
    LocalMux I__4580 (
            .O(N__18961),
            .I(N__18946));
    InMux I__4579 (
            .O(N__18960),
            .I(N__18943));
    InMux I__4578 (
            .O(N__18959),
            .I(N__18938));
    InMux I__4577 (
            .O(N__18956),
            .I(N__18938));
    InMux I__4576 (
            .O(N__18955),
            .I(N__18933));
    InMux I__4575 (
            .O(N__18954),
            .I(N__18933));
    InMux I__4574 (
            .O(N__18953),
            .I(N__18928));
    InMux I__4573 (
            .O(N__18952),
            .I(N__18928));
    Span4Mux_h I__4572 (
            .O(N__18949),
            .I(N__18925));
    Span4Mux_h I__4571 (
            .O(N__18946),
            .I(N__18918));
    LocalMux I__4570 (
            .O(N__18943),
            .I(N__18918));
    LocalMux I__4569 (
            .O(N__18938),
            .I(N__18918));
    LocalMux I__4568 (
            .O(N__18933),
            .I(\Lab_UT.state_i_3_2 ));
    LocalMux I__4567 (
            .O(N__18928),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4566 (
            .O(N__18925),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4565 (
            .O(N__18918),
            .I(\Lab_UT.state_i_3_2 ));
    InMux I__4564 (
            .O(N__18909),
            .I(N__18905));
    InMux I__4563 (
            .O(N__18908),
            .I(N__18897));
    LocalMux I__4562 (
            .O(N__18905),
            .I(N__18890));
    InMux I__4561 (
            .O(N__18904),
            .I(N__18887));
    InMux I__4560 (
            .O(N__18903),
            .I(N__18878));
    InMux I__4559 (
            .O(N__18902),
            .I(N__18878));
    InMux I__4558 (
            .O(N__18901),
            .I(N__18878));
    InMux I__4557 (
            .O(N__18900),
            .I(N__18878));
    LocalMux I__4556 (
            .O(N__18897),
            .I(N__18874));
    InMux I__4555 (
            .O(N__18896),
            .I(N__18865));
    InMux I__4554 (
            .O(N__18895),
            .I(N__18865));
    InMux I__4553 (
            .O(N__18894),
            .I(N__18865));
    InMux I__4552 (
            .O(N__18893),
            .I(N__18865));
    Span4Mux_h I__4551 (
            .O(N__18890),
            .I(N__18858));
    LocalMux I__4550 (
            .O(N__18887),
            .I(N__18858));
    LocalMux I__4549 (
            .O(N__18878),
            .I(N__18858));
    InMux I__4548 (
            .O(N__18877),
            .I(N__18855));
    Odrv4 I__4547 (
            .O(N__18874),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4546 (
            .O(N__18865),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__4545 (
            .O(N__18858),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4544 (
            .O(N__18855),
            .I(\Lab_UT.state_0 ));
    InMux I__4543 (
            .O(N__18846),
            .I(N__18836));
    InMux I__4542 (
            .O(N__18845),
            .I(N__18836));
    InMux I__4541 (
            .O(N__18844),
            .I(N__18836));
    InMux I__4540 (
            .O(N__18843),
            .I(N__18833));
    LocalMux I__4539 (
            .O(N__18836),
            .I(N__18830));
    LocalMux I__4538 (
            .O(N__18833),
            .I(N__18827));
    Odrv4 I__4537 (
            .O(N__18830),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    Odrv4 I__4536 (
            .O(N__18827),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__4535 (
            .O(N__18822),
            .I(N__18819));
    LocalMux I__4534 (
            .O(N__18819),
            .I(N__18816));
    Span4Mux_h I__4533 (
            .O(N__18816),
            .I(N__18811));
    InMux I__4532 (
            .O(N__18815),
            .I(N__18808));
    InMux I__4531 (
            .O(N__18814),
            .I(N__18805));
    Odrv4 I__4530 (
            .O(N__18811),
            .I(\Lab_UT.nine ));
    LocalMux I__4529 (
            .O(N__18808),
            .I(\Lab_UT.nine ));
    LocalMux I__4528 (
            .O(N__18805),
            .I(\Lab_UT.nine ));
    InMux I__4527 (
            .O(N__18798),
            .I(N__18788));
    InMux I__4526 (
            .O(N__18797),
            .I(N__18788));
    InMux I__4525 (
            .O(N__18796),
            .I(N__18788));
    InMux I__4524 (
            .O(N__18795),
            .I(N__18785));
    LocalMux I__4523 (
            .O(N__18788),
            .I(N__18782));
    LocalMux I__4522 (
            .O(N__18785),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    Odrv4 I__4521 (
            .O(N__18782),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    InMux I__4520 (
            .O(N__18777),
            .I(N__18772));
    InMux I__4519 (
            .O(N__18776),
            .I(N__18767));
    InMux I__4518 (
            .O(N__18775),
            .I(N__18767));
    LocalMux I__4517 (
            .O(N__18772),
            .I(N__18761));
    LocalMux I__4516 (
            .O(N__18767),
            .I(N__18761));
    InMux I__4515 (
            .O(N__18766),
            .I(N__18758));
    Span4Mux_h I__4514 (
            .O(N__18761),
            .I(N__18755));
    LocalMux I__4513 (
            .O(N__18758),
            .I(\Lab_UT.q_RNI84NN1_2 ));
    Odrv4 I__4512 (
            .O(N__18755),
            .I(\Lab_UT.q_RNI84NN1_2 ));
    InMux I__4511 (
            .O(N__18750),
            .I(N__18738));
    InMux I__4510 (
            .O(N__18749),
            .I(N__18735));
    InMux I__4509 (
            .O(N__18748),
            .I(N__18732));
    InMux I__4508 (
            .O(N__18747),
            .I(N__18729));
    InMux I__4507 (
            .O(N__18746),
            .I(N__18726));
    InMux I__4506 (
            .O(N__18745),
            .I(N__18719));
    InMux I__4505 (
            .O(N__18744),
            .I(N__18719));
    InMux I__4504 (
            .O(N__18743),
            .I(N__18719));
    SRMux I__4503 (
            .O(N__18742),
            .I(N__18714));
    InMux I__4502 (
            .O(N__18741),
            .I(N__18714));
    LocalMux I__4501 (
            .O(N__18738),
            .I(N__18684));
    LocalMux I__4500 (
            .O(N__18735),
            .I(N__18681));
    LocalMux I__4499 (
            .O(N__18732),
            .I(N__18678));
    LocalMux I__4498 (
            .O(N__18729),
            .I(N__18675));
    LocalMux I__4497 (
            .O(N__18726),
            .I(N__18672));
    LocalMux I__4496 (
            .O(N__18719),
            .I(N__18669));
    LocalMux I__4495 (
            .O(N__18714),
            .I(N__18645));
    SRMux I__4494 (
            .O(N__18713),
            .I(N__18534));
    SRMux I__4493 (
            .O(N__18712),
            .I(N__18534));
    SRMux I__4492 (
            .O(N__18711),
            .I(N__18534));
    SRMux I__4491 (
            .O(N__18710),
            .I(N__18534));
    SRMux I__4490 (
            .O(N__18709),
            .I(N__18534));
    SRMux I__4489 (
            .O(N__18708),
            .I(N__18534));
    SRMux I__4488 (
            .O(N__18707),
            .I(N__18534));
    SRMux I__4487 (
            .O(N__18706),
            .I(N__18534));
    SRMux I__4486 (
            .O(N__18705),
            .I(N__18534));
    SRMux I__4485 (
            .O(N__18704),
            .I(N__18534));
    SRMux I__4484 (
            .O(N__18703),
            .I(N__18534));
    SRMux I__4483 (
            .O(N__18702),
            .I(N__18534));
    SRMux I__4482 (
            .O(N__18701),
            .I(N__18534));
    SRMux I__4481 (
            .O(N__18700),
            .I(N__18534));
    SRMux I__4480 (
            .O(N__18699),
            .I(N__18534));
    SRMux I__4479 (
            .O(N__18698),
            .I(N__18534));
    SRMux I__4478 (
            .O(N__18697),
            .I(N__18534));
    SRMux I__4477 (
            .O(N__18696),
            .I(N__18534));
    SRMux I__4476 (
            .O(N__18695),
            .I(N__18534));
    SRMux I__4475 (
            .O(N__18694),
            .I(N__18534));
    SRMux I__4474 (
            .O(N__18693),
            .I(N__18534));
    SRMux I__4473 (
            .O(N__18692),
            .I(N__18534));
    SRMux I__4472 (
            .O(N__18691),
            .I(N__18534));
    SRMux I__4471 (
            .O(N__18690),
            .I(N__18534));
    SRMux I__4470 (
            .O(N__18689),
            .I(N__18534));
    SRMux I__4469 (
            .O(N__18688),
            .I(N__18534));
    SRMux I__4468 (
            .O(N__18687),
            .I(N__18534));
    Glb2LocalMux I__4467 (
            .O(N__18684),
            .I(N__18534));
    Glb2LocalMux I__4466 (
            .O(N__18681),
            .I(N__18534));
    Glb2LocalMux I__4465 (
            .O(N__18678),
            .I(N__18534));
    Glb2LocalMux I__4464 (
            .O(N__18675),
            .I(N__18534));
    Glb2LocalMux I__4463 (
            .O(N__18672),
            .I(N__18534));
    Glb2LocalMux I__4462 (
            .O(N__18669),
            .I(N__18534));
    SRMux I__4461 (
            .O(N__18668),
            .I(N__18534));
    SRMux I__4460 (
            .O(N__18667),
            .I(N__18534));
    SRMux I__4459 (
            .O(N__18666),
            .I(N__18534));
    SRMux I__4458 (
            .O(N__18665),
            .I(N__18534));
    SRMux I__4457 (
            .O(N__18664),
            .I(N__18534));
    SRMux I__4456 (
            .O(N__18663),
            .I(N__18534));
    SRMux I__4455 (
            .O(N__18662),
            .I(N__18534));
    SRMux I__4454 (
            .O(N__18661),
            .I(N__18534));
    SRMux I__4453 (
            .O(N__18660),
            .I(N__18534));
    SRMux I__4452 (
            .O(N__18659),
            .I(N__18534));
    SRMux I__4451 (
            .O(N__18658),
            .I(N__18534));
    SRMux I__4450 (
            .O(N__18657),
            .I(N__18534));
    SRMux I__4449 (
            .O(N__18656),
            .I(N__18534));
    SRMux I__4448 (
            .O(N__18655),
            .I(N__18534));
    SRMux I__4447 (
            .O(N__18654),
            .I(N__18534));
    SRMux I__4446 (
            .O(N__18653),
            .I(N__18534));
    SRMux I__4445 (
            .O(N__18652),
            .I(N__18534));
    SRMux I__4444 (
            .O(N__18651),
            .I(N__18534));
    SRMux I__4443 (
            .O(N__18650),
            .I(N__18534));
    SRMux I__4442 (
            .O(N__18649),
            .I(N__18534));
    SRMux I__4441 (
            .O(N__18648),
            .I(N__18534));
    Glb2LocalMux I__4440 (
            .O(N__18645),
            .I(N__18534));
    GlobalMux I__4439 (
            .O(N__18534),
            .I(N__18531));
    gio2CtrlBuf I__4438 (
            .O(N__18531),
            .I(rst_g));
    CascadeMux I__4437 (
            .O(N__18528),
            .I(N__18523));
    InMux I__4436 (
            .O(N__18527),
            .I(N__18517));
    InMux I__4435 (
            .O(N__18526),
            .I(N__18517));
    InMux I__4434 (
            .O(N__18523),
            .I(N__18512));
    InMux I__4433 (
            .O(N__18522),
            .I(N__18512));
    LocalMux I__4432 (
            .O(N__18517),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    LocalMux I__4431 (
            .O(N__18512),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    ClkMux I__4430 (
            .O(N__18507),
            .I(N__18252));
    ClkMux I__4429 (
            .O(N__18506),
            .I(N__18252));
    ClkMux I__4428 (
            .O(N__18505),
            .I(N__18252));
    ClkMux I__4427 (
            .O(N__18504),
            .I(N__18252));
    ClkMux I__4426 (
            .O(N__18503),
            .I(N__18252));
    ClkMux I__4425 (
            .O(N__18502),
            .I(N__18252));
    ClkMux I__4424 (
            .O(N__18501),
            .I(N__18252));
    ClkMux I__4423 (
            .O(N__18500),
            .I(N__18252));
    ClkMux I__4422 (
            .O(N__18499),
            .I(N__18252));
    ClkMux I__4421 (
            .O(N__18498),
            .I(N__18252));
    ClkMux I__4420 (
            .O(N__18497),
            .I(N__18252));
    ClkMux I__4419 (
            .O(N__18496),
            .I(N__18252));
    ClkMux I__4418 (
            .O(N__18495),
            .I(N__18252));
    ClkMux I__4417 (
            .O(N__18494),
            .I(N__18252));
    ClkMux I__4416 (
            .O(N__18493),
            .I(N__18252));
    ClkMux I__4415 (
            .O(N__18492),
            .I(N__18252));
    ClkMux I__4414 (
            .O(N__18491),
            .I(N__18252));
    ClkMux I__4413 (
            .O(N__18490),
            .I(N__18252));
    ClkMux I__4412 (
            .O(N__18489),
            .I(N__18252));
    ClkMux I__4411 (
            .O(N__18488),
            .I(N__18252));
    ClkMux I__4410 (
            .O(N__18487),
            .I(N__18252));
    ClkMux I__4409 (
            .O(N__18486),
            .I(N__18252));
    ClkMux I__4408 (
            .O(N__18485),
            .I(N__18252));
    ClkMux I__4407 (
            .O(N__18484),
            .I(N__18252));
    ClkMux I__4406 (
            .O(N__18483),
            .I(N__18252));
    ClkMux I__4405 (
            .O(N__18482),
            .I(N__18252));
    ClkMux I__4404 (
            .O(N__18481),
            .I(N__18252));
    ClkMux I__4403 (
            .O(N__18480),
            .I(N__18252));
    ClkMux I__4402 (
            .O(N__18479),
            .I(N__18252));
    ClkMux I__4401 (
            .O(N__18478),
            .I(N__18252));
    ClkMux I__4400 (
            .O(N__18477),
            .I(N__18252));
    ClkMux I__4399 (
            .O(N__18476),
            .I(N__18252));
    ClkMux I__4398 (
            .O(N__18475),
            .I(N__18252));
    ClkMux I__4397 (
            .O(N__18474),
            .I(N__18252));
    ClkMux I__4396 (
            .O(N__18473),
            .I(N__18252));
    ClkMux I__4395 (
            .O(N__18472),
            .I(N__18252));
    ClkMux I__4394 (
            .O(N__18471),
            .I(N__18252));
    ClkMux I__4393 (
            .O(N__18470),
            .I(N__18252));
    ClkMux I__4392 (
            .O(N__18469),
            .I(N__18252));
    ClkMux I__4391 (
            .O(N__18468),
            .I(N__18252));
    ClkMux I__4390 (
            .O(N__18467),
            .I(N__18252));
    ClkMux I__4389 (
            .O(N__18466),
            .I(N__18252));
    ClkMux I__4388 (
            .O(N__18465),
            .I(N__18252));
    ClkMux I__4387 (
            .O(N__18464),
            .I(N__18252));
    ClkMux I__4386 (
            .O(N__18463),
            .I(N__18252));
    ClkMux I__4385 (
            .O(N__18462),
            .I(N__18252));
    ClkMux I__4384 (
            .O(N__18461),
            .I(N__18252));
    ClkMux I__4383 (
            .O(N__18460),
            .I(N__18252));
    ClkMux I__4382 (
            .O(N__18459),
            .I(N__18252));
    ClkMux I__4381 (
            .O(N__18458),
            .I(N__18252));
    ClkMux I__4380 (
            .O(N__18457),
            .I(N__18252));
    ClkMux I__4379 (
            .O(N__18456),
            .I(N__18252));
    ClkMux I__4378 (
            .O(N__18455),
            .I(N__18252));
    ClkMux I__4377 (
            .O(N__18454),
            .I(N__18252));
    ClkMux I__4376 (
            .O(N__18453),
            .I(N__18252));
    ClkMux I__4375 (
            .O(N__18452),
            .I(N__18252));
    ClkMux I__4374 (
            .O(N__18451),
            .I(N__18252));
    ClkMux I__4373 (
            .O(N__18450),
            .I(N__18252));
    ClkMux I__4372 (
            .O(N__18449),
            .I(N__18252));
    ClkMux I__4371 (
            .O(N__18448),
            .I(N__18252));
    ClkMux I__4370 (
            .O(N__18447),
            .I(N__18252));
    ClkMux I__4369 (
            .O(N__18446),
            .I(N__18252));
    ClkMux I__4368 (
            .O(N__18445),
            .I(N__18252));
    ClkMux I__4367 (
            .O(N__18444),
            .I(N__18252));
    ClkMux I__4366 (
            .O(N__18443),
            .I(N__18252));
    ClkMux I__4365 (
            .O(N__18442),
            .I(N__18252));
    ClkMux I__4364 (
            .O(N__18441),
            .I(N__18252));
    ClkMux I__4363 (
            .O(N__18440),
            .I(N__18252));
    ClkMux I__4362 (
            .O(N__18439),
            .I(N__18252));
    ClkMux I__4361 (
            .O(N__18438),
            .I(N__18252));
    ClkMux I__4360 (
            .O(N__18437),
            .I(N__18252));
    ClkMux I__4359 (
            .O(N__18436),
            .I(N__18252));
    ClkMux I__4358 (
            .O(N__18435),
            .I(N__18252));
    ClkMux I__4357 (
            .O(N__18434),
            .I(N__18252));
    ClkMux I__4356 (
            .O(N__18433),
            .I(N__18252));
    ClkMux I__4355 (
            .O(N__18432),
            .I(N__18252));
    ClkMux I__4354 (
            .O(N__18431),
            .I(N__18252));
    ClkMux I__4353 (
            .O(N__18430),
            .I(N__18252));
    ClkMux I__4352 (
            .O(N__18429),
            .I(N__18252));
    ClkMux I__4351 (
            .O(N__18428),
            .I(N__18252));
    ClkMux I__4350 (
            .O(N__18427),
            .I(N__18252));
    ClkMux I__4349 (
            .O(N__18426),
            .I(N__18252));
    ClkMux I__4348 (
            .O(N__18425),
            .I(N__18252));
    ClkMux I__4347 (
            .O(N__18424),
            .I(N__18252));
    ClkMux I__4346 (
            .O(N__18423),
            .I(N__18252));
    GlobalMux I__4345 (
            .O(N__18252),
            .I(N__18249));
    gio2CtrlBuf I__4344 (
            .O(N__18249),
            .I(clk_g));
    SRMux I__4343 (
            .O(N__18246),
            .I(N__18243));
    LocalMux I__4342 (
            .O(N__18243),
            .I(N__18239));
    SRMux I__4341 (
            .O(N__18242),
            .I(N__18236));
    Span4Mux_v I__4340 (
            .O(N__18239),
            .I(N__18230));
    LocalMux I__4339 (
            .O(N__18236),
            .I(N__18230));
    SRMux I__4338 (
            .O(N__18235),
            .I(N__18227));
    Span4Mux_v I__4337 (
            .O(N__18230),
            .I(N__18224));
    LocalMux I__4336 (
            .O(N__18227),
            .I(N__18220));
    IoSpan4Mux I__4335 (
            .O(N__18224),
            .I(N__18217));
    SRMux I__4334 (
            .O(N__18223),
            .I(N__18214));
    Span4Mux_v I__4333 (
            .O(N__18220),
            .I(N__18211));
    Span4Mux_s2_h I__4332 (
            .O(N__18217),
            .I(N__18206));
    LocalMux I__4331 (
            .O(N__18214),
            .I(N__18206));
    Span4Mux_h I__4330 (
            .O(N__18211),
            .I(N__18201));
    Span4Mux_h I__4329 (
            .O(N__18206),
            .I(N__18201));
    Span4Mux_h I__4328 (
            .O(N__18201),
            .I(N__18198));
    Odrv4 I__4327 (
            .O(N__18198),
            .I(oneSecStrb_i));
    InMux I__4326 (
            .O(N__18195),
            .I(N__18192));
    LocalMux I__4325 (
            .O(N__18192),
            .I(N__18189));
    Span4Mux_h I__4324 (
            .O(N__18189),
            .I(N__18186));
    Odrv4 I__4323 (
            .O(N__18186),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_4 ));
    CascadeMux I__4322 (
            .O(N__18183),
            .I(\Lab_UT.three_2_cascade_ ));
    InMux I__4321 (
            .O(N__18180),
            .I(N__18175));
    CascadeMux I__4320 (
            .O(N__18179),
            .I(N__18172));
    CascadeMux I__4319 (
            .O(N__18178),
            .I(N__18167));
    LocalMux I__4318 (
            .O(N__18175),
            .I(N__18163));
    InMux I__4317 (
            .O(N__18172),
            .I(N__18150));
    InMux I__4316 (
            .O(N__18171),
            .I(N__18150));
    InMux I__4315 (
            .O(N__18170),
            .I(N__18150));
    InMux I__4314 (
            .O(N__18167),
            .I(N__18145));
    InMux I__4313 (
            .O(N__18166),
            .I(N__18145));
    Span4Mux_h I__4312 (
            .O(N__18163),
            .I(N__18142));
    InMux I__4311 (
            .O(N__18162),
            .I(N__18137));
    InMux I__4310 (
            .O(N__18161),
            .I(N__18137));
    InMux I__4309 (
            .O(N__18160),
            .I(N__18130));
    InMux I__4308 (
            .O(N__18159),
            .I(N__18130));
    InMux I__4307 (
            .O(N__18158),
            .I(N__18130));
    InMux I__4306 (
            .O(N__18157),
            .I(N__18127));
    LocalMux I__4305 (
            .O(N__18150),
            .I(N__18122));
    LocalMux I__4304 (
            .O(N__18145),
            .I(N__18122));
    Odrv4 I__4303 (
            .O(N__18142),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__4302 (
            .O(N__18137),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__4301 (
            .O(N__18130),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__4300 (
            .O(N__18127),
            .I(\Lab_UT.di_Stens_1 ));
    Odrv12 I__4299 (
            .O(N__18122),
            .I(\Lab_UT.di_Stens_1 ));
    CascadeMux I__4298 (
            .O(N__18111),
            .I(N__18108));
    InMux I__4297 (
            .O(N__18108),
            .I(N__18105));
    LocalMux I__4296 (
            .O(N__18105),
            .I(N__18102));
    Odrv4 I__4295 (
            .O(N__18102),
            .I(\Lab_UT.didp.countrce2.un15_ce_2 ));
    CascadeMux I__4294 (
            .O(N__18099),
            .I(\Lab_UT.didp.countrce2.un15_ce_2_cascade_ ));
    InMux I__4293 (
            .O(N__18096),
            .I(N__18092));
    InMux I__4292 (
            .O(N__18095),
            .I(N__18077));
    LocalMux I__4291 (
            .O(N__18092),
            .I(N__18074));
    InMux I__4290 (
            .O(N__18091),
            .I(N__18069));
    InMux I__4289 (
            .O(N__18090),
            .I(N__18069));
    InMux I__4288 (
            .O(N__18089),
            .I(N__18062));
    InMux I__4287 (
            .O(N__18088),
            .I(N__18062));
    InMux I__4286 (
            .O(N__18087),
            .I(N__18062));
    InMux I__4285 (
            .O(N__18086),
            .I(N__18055));
    InMux I__4284 (
            .O(N__18085),
            .I(N__18055));
    InMux I__4283 (
            .O(N__18084),
            .I(N__18055));
    InMux I__4282 (
            .O(N__18083),
            .I(N__18046));
    InMux I__4281 (
            .O(N__18082),
            .I(N__18046));
    InMux I__4280 (
            .O(N__18081),
            .I(N__18046));
    InMux I__4279 (
            .O(N__18080),
            .I(N__18046));
    LocalMux I__4278 (
            .O(N__18077),
            .I(N__18037));
    Span12Mux_s6_h I__4277 (
            .O(N__18074),
            .I(N__18037));
    LocalMux I__4276 (
            .O(N__18069),
            .I(N__18037));
    LocalMux I__4275 (
            .O(N__18062),
            .I(N__18037));
    LocalMux I__4274 (
            .O(N__18055),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__4273 (
            .O(N__18046),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv12 I__4272 (
            .O(N__18037),
            .I(\Lab_UT.di_Stens_0 ));
    CascadeMux I__4271 (
            .O(N__18030),
            .I(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ));
    CascadeMux I__4270 (
            .O(N__18027),
            .I(N__18022));
    InMux I__4269 (
            .O(N__18026),
            .I(N__18012));
    InMux I__4268 (
            .O(N__18025),
            .I(N__18007));
    InMux I__4267 (
            .O(N__18022),
            .I(N__18007));
    CascadeMux I__4266 (
            .O(N__18021),
            .I(N__18004));
    CascadeMux I__4265 (
            .O(N__18020),
            .I(N__18000));
    CascadeMux I__4264 (
            .O(N__18019),
            .I(N__17997));
    CascadeMux I__4263 (
            .O(N__18018),
            .I(N__17994));
    CascadeMux I__4262 (
            .O(N__18017),
            .I(N__17991));
    InMux I__4261 (
            .O(N__18016),
            .I(N__17986));
    InMux I__4260 (
            .O(N__18015),
            .I(N__17986));
    LocalMux I__4259 (
            .O(N__18012),
            .I(N__17981));
    LocalMux I__4258 (
            .O(N__18007),
            .I(N__17981));
    InMux I__4257 (
            .O(N__18004),
            .I(N__17974));
    InMux I__4256 (
            .O(N__18003),
            .I(N__17974));
    InMux I__4255 (
            .O(N__18000),
            .I(N__17974));
    InMux I__4254 (
            .O(N__17997),
            .I(N__17971));
    InMux I__4253 (
            .O(N__17994),
            .I(N__17966));
    InMux I__4252 (
            .O(N__17991),
            .I(N__17966));
    LocalMux I__4251 (
            .O(N__17986),
            .I(N__17961));
    Span4Mux_h I__4250 (
            .O(N__17981),
            .I(N__17961));
    LocalMux I__4249 (
            .O(N__17974),
            .I(N__17958));
    LocalMux I__4248 (
            .O(N__17971),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4247 (
            .O(N__17966),
            .I(\Lab_UT.di_Stens_3 ));
    Odrv4 I__4246 (
            .O(N__17961),
            .I(\Lab_UT.di_Stens_3 ));
    Odrv12 I__4245 (
            .O(N__17958),
            .I(\Lab_UT.di_Stens_3 ));
    InMux I__4244 (
            .O(N__17949),
            .I(N__17940));
    InMux I__4243 (
            .O(N__17948),
            .I(N__17940));
    InMux I__4242 (
            .O(N__17947),
            .I(N__17937));
    InMux I__4241 (
            .O(N__17946),
            .I(N__17934));
    InMux I__4240 (
            .O(N__17945),
            .I(N__17931));
    LocalMux I__4239 (
            .O(N__17940),
            .I(N__17928));
    LocalMux I__4238 (
            .O(N__17937),
            .I(\Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ));
    LocalMux I__4237 (
            .O(N__17934),
            .I(\Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ));
    LocalMux I__4236 (
            .O(N__17931),
            .I(\Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ));
    Odrv4 I__4235 (
            .O(N__17928),
            .I(\Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ));
    InMux I__4234 (
            .O(N__17919),
            .I(N__17916));
    LocalMux I__4233 (
            .O(N__17916),
            .I(N__17913));
    Span4Mux_h I__4232 (
            .O(N__17913),
            .I(N__17908));
    InMux I__4231 (
            .O(N__17912),
            .I(N__17905));
    InMux I__4230 (
            .O(N__17911),
            .I(N__17902));
    Odrv4 I__4229 (
            .O(N__17908),
            .I(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1 ));
    LocalMux I__4228 (
            .O(N__17905),
            .I(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1 ));
    LocalMux I__4227 (
            .O(N__17902),
            .I(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1 ));
    CascadeMux I__4226 (
            .O(N__17895),
            .I(N__17891));
    CascadeMux I__4225 (
            .O(N__17894),
            .I(N__17888));
    InMux I__4224 (
            .O(N__17891),
            .I(N__17881));
    InMux I__4223 (
            .O(N__17888),
            .I(N__17881));
    InMux I__4222 (
            .O(N__17887),
            .I(N__17878));
    CascadeMux I__4221 (
            .O(N__17886),
            .I(N__17871));
    LocalMux I__4220 (
            .O(N__17881),
            .I(N__17865));
    LocalMux I__4219 (
            .O(N__17878),
            .I(N__17865));
    InMux I__4218 (
            .O(N__17877),
            .I(N__17862));
    CascadeMux I__4217 (
            .O(N__17876),
            .I(N__17856));
    InMux I__4216 (
            .O(N__17875),
            .I(N__17849));
    InMux I__4215 (
            .O(N__17874),
            .I(N__17849));
    InMux I__4214 (
            .O(N__17871),
            .I(N__17849));
    CascadeMux I__4213 (
            .O(N__17870),
            .I(N__17846));
    Span4Mux_v I__4212 (
            .O(N__17865),
            .I(N__17841));
    LocalMux I__4211 (
            .O(N__17862),
            .I(N__17841));
    InMux I__4210 (
            .O(N__17861),
            .I(N__17832));
    InMux I__4209 (
            .O(N__17860),
            .I(N__17832));
    InMux I__4208 (
            .O(N__17859),
            .I(N__17832));
    InMux I__4207 (
            .O(N__17856),
            .I(N__17832));
    LocalMux I__4206 (
            .O(N__17849),
            .I(N__17829));
    InMux I__4205 (
            .O(N__17846),
            .I(N__17826));
    Span4Mux_h I__4204 (
            .O(N__17841),
            .I(N__17823));
    LocalMux I__4203 (
            .O(N__17832),
            .I(N__17816));
    Span4Mux_v I__4202 (
            .O(N__17829),
            .I(N__17816));
    LocalMux I__4201 (
            .O(N__17826),
            .I(N__17816));
    Sp12to4 I__4200 (
            .O(N__17823),
            .I(N__17813));
    Span4Mux_h I__4199 (
            .O(N__17816),
            .I(N__17810));
    Odrv12 I__4198 (
            .O(N__17813),
            .I(\Lab_UT.dictrl.state_retZ0Z_4 ));
    Odrv4 I__4197 (
            .O(N__17810),
            .I(\Lab_UT.dictrl.state_retZ0Z_4 ));
    InMux I__4196 (
            .O(N__17805),
            .I(N__17800));
    InMux I__4195 (
            .O(N__17804),
            .I(N__17797));
    InMux I__4194 (
            .O(N__17803),
            .I(N__17793));
    LocalMux I__4193 (
            .O(N__17800),
            .I(N__17790));
    LocalMux I__4192 (
            .O(N__17797),
            .I(N__17787));
    InMux I__4191 (
            .O(N__17796),
            .I(N__17784));
    LocalMux I__4190 (
            .O(N__17793),
            .I(\Lab_UT.dictrl.next_state_set_0 ));
    Odrv4 I__4189 (
            .O(N__17790),
            .I(\Lab_UT.dictrl.next_state_set_0 ));
    Odrv4 I__4188 (
            .O(N__17787),
            .I(\Lab_UT.dictrl.next_state_set_0 ));
    LocalMux I__4187 (
            .O(N__17784),
            .I(\Lab_UT.dictrl.next_state_set_0 ));
    InMux I__4186 (
            .O(N__17775),
            .I(N__17770));
    InMux I__4185 (
            .O(N__17774),
            .I(N__17765));
    InMux I__4184 (
            .O(N__17773),
            .I(N__17765));
    LocalMux I__4183 (
            .O(N__17770),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__4182 (
            .O(N__17765),
            .I(\Lab_UT.state_i_3_1 ));
    CascadeMux I__4181 (
            .O(N__17760),
            .I(N__17757));
    InMux I__4180 (
            .O(N__17757),
            .I(N__17753));
    InMux I__4179 (
            .O(N__17756),
            .I(N__17749));
    LocalMux I__4178 (
            .O(N__17753),
            .I(N__17746));
    InMux I__4177 (
            .O(N__17752),
            .I(N__17743));
    LocalMux I__4176 (
            .O(N__17749),
            .I(N__17736));
    Span4Mux_v I__4175 (
            .O(N__17746),
            .I(N__17731));
    LocalMux I__4174 (
            .O(N__17743),
            .I(N__17731));
    InMux I__4173 (
            .O(N__17742),
            .I(N__17726));
    InMux I__4172 (
            .O(N__17741),
            .I(N__17726));
    InMux I__4171 (
            .O(N__17740),
            .I(N__17723));
    InMux I__4170 (
            .O(N__17739),
            .I(N__17720));
    Odrv4 I__4169 (
            .O(N__17736),
            .I(bu_rx_data_3));
    Odrv4 I__4168 (
            .O(N__17731),
            .I(bu_rx_data_3));
    LocalMux I__4167 (
            .O(N__17726),
            .I(bu_rx_data_3));
    LocalMux I__4166 (
            .O(N__17723),
            .I(bu_rx_data_3));
    LocalMux I__4165 (
            .O(N__17720),
            .I(bu_rx_data_3));
    InMux I__4164 (
            .O(N__17709),
            .I(N__17705));
    InMux I__4163 (
            .O(N__17708),
            .I(N__17698));
    LocalMux I__4162 (
            .O(N__17705),
            .I(N__17695));
    InMux I__4161 (
            .O(N__17704),
            .I(N__17692));
    InMux I__4160 (
            .O(N__17703),
            .I(N__17687));
    InMux I__4159 (
            .O(N__17702),
            .I(N__17687));
    CascadeMux I__4158 (
            .O(N__17701),
            .I(N__17683));
    LocalMux I__4157 (
            .O(N__17698),
            .I(N__17674));
    Span4Mux_h I__4156 (
            .O(N__17695),
            .I(N__17674));
    LocalMux I__4155 (
            .O(N__17692),
            .I(N__17674));
    LocalMux I__4154 (
            .O(N__17687),
            .I(N__17674));
    InMux I__4153 (
            .O(N__17686),
            .I(N__17669));
    InMux I__4152 (
            .O(N__17683),
            .I(N__17669));
    Span4Mux_v I__4151 (
            .O(N__17674),
            .I(N__17664));
    LocalMux I__4150 (
            .O(N__17669),
            .I(N__17664));
    Odrv4 I__4149 (
            .O(N__17664),
            .I(bu_rx_data_2));
    CEMux I__4148 (
            .O(N__17661),
            .I(N__17657));
    CEMux I__4147 (
            .O(N__17660),
            .I(N__17654));
    LocalMux I__4146 (
            .O(N__17657),
            .I(N__17649));
    LocalMux I__4145 (
            .O(N__17654),
            .I(N__17646));
    CEMux I__4144 (
            .O(N__17653),
            .I(N__17643));
    CEMux I__4143 (
            .O(N__17652),
            .I(N__17640));
    Span4Mux_v I__4142 (
            .O(N__17649),
            .I(N__17637));
    Span4Mux_v I__4141 (
            .O(N__17646),
            .I(N__17634));
    LocalMux I__4140 (
            .O(N__17643),
            .I(N__17631));
    LocalMux I__4139 (
            .O(N__17640),
            .I(N__17628));
    Span4Mux_h I__4138 (
            .O(N__17637),
            .I(N__17625));
    Span4Mux_h I__4137 (
            .O(N__17634),
            .I(N__17622));
    Span4Mux_h I__4136 (
            .O(N__17631),
            .I(N__17619));
    Span4Mux_v I__4135 (
            .O(N__17628),
            .I(N__17616));
    Odrv4 I__4134 (
            .O(N__17625),
            .I(\buart.Z_rx.sample ));
    Odrv4 I__4133 (
            .O(N__17622),
            .I(\buart.Z_rx.sample ));
    Odrv4 I__4132 (
            .O(N__17619),
            .I(\buart.Z_rx.sample ));
    Odrv4 I__4131 (
            .O(N__17616),
            .I(\buart.Z_rx.sample ));
    InMux I__4130 (
            .O(N__17607),
            .I(N__17604));
    LocalMux I__4129 (
            .O(N__17604),
            .I(N__17601));
    Odrv4 I__4128 (
            .O(N__17601),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_0 ));
    InMux I__4127 (
            .O(N__17598),
            .I(N__17595));
    LocalMux I__4126 (
            .O(N__17595),
            .I(N__17592));
    Odrv4 I__4125 (
            .O(N__17592),
            .I(\Lab_UT.bcd2segment1.N_192 ));
    InMux I__4124 (
            .O(N__17589),
            .I(N__17586));
    LocalMux I__4123 (
            .O(N__17586),
            .I(N__17583));
    Span4Mux_s3_v I__4122 (
            .O(N__17583),
            .I(N__17580));
    Span4Mux_v I__4121 (
            .O(N__17580),
            .I(N__17577));
    Odrv4 I__4120 (
            .O(N__17577),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_5 ));
    InMux I__4119 (
            .O(N__17574),
            .I(N__17571));
    LocalMux I__4118 (
            .O(N__17571),
            .I(N__17568));
    Odrv4 I__4117 (
            .O(N__17568),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_3 ));
    CascadeMux I__4116 (
            .O(N__17565),
            .I(N__17562));
    InMux I__4115 (
            .O(N__17562),
            .I(N__17558));
    CascadeMux I__4114 (
            .O(N__17561),
            .I(N__17555));
    LocalMux I__4113 (
            .O(N__17558),
            .I(N__17552));
    InMux I__4112 (
            .O(N__17555),
            .I(N__17549));
    Span4Mux_v I__4111 (
            .O(N__17552),
            .I(N__17542));
    LocalMux I__4110 (
            .O(N__17549),
            .I(N__17542));
    InMux I__4109 (
            .O(N__17548),
            .I(N__17539));
    InMux I__4108 (
            .O(N__17547),
            .I(N__17536));
    Odrv4 I__4107 (
            .O(N__17542),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    LocalMux I__4106 (
            .O(N__17539),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    LocalMux I__4105 (
            .O(N__17536),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    InMux I__4104 (
            .O(N__17529),
            .I(N__17526));
    LocalMux I__4103 (
            .O(N__17526),
            .I(N__17522));
    InMux I__4102 (
            .O(N__17525),
            .I(N__17517));
    Span4Mux_h I__4101 (
            .O(N__17522),
            .I(N__17514));
    InMux I__4100 (
            .O(N__17521),
            .I(N__17511));
    InMux I__4099 (
            .O(N__17520),
            .I(N__17508));
    LocalMux I__4098 (
            .O(N__17517),
            .I(N__17505));
    Odrv4 I__4097 (
            .O(N__17514),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    LocalMux I__4096 (
            .O(N__17511),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    LocalMux I__4095 (
            .O(N__17508),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    Odrv4 I__4094 (
            .O(N__17505),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    CEMux I__4093 (
            .O(N__17496),
            .I(N__17490));
    CEMux I__4092 (
            .O(N__17495),
            .I(N__17487));
    CEMux I__4091 (
            .O(N__17494),
            .I(N__17484));
    CEMux I__4090 (
            .O(N__17493),
            .I(N__17481));
    LocalMux I__4089 (
            .O(N__17490),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    LocalMux I__4088 (
            .O(N__17487),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    LocalMux I__4087 (
            .O(N__17484),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    LocalMux I__4086 (
            .O(N__17481),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    SRMux I__4085 (
            .O(N__17472),
            .I(N__17469));
    LocalMux I__4084 (
            .O(N__17469),
            .I(N__17466));
    Span4Mux_h I__4083 (
            .O(N__17466),
            .I(N__17462));
    InMux I__4082 (
            .O(N__17465),
            .I(N__17459));
    Odrv4 I__4081 (
            .O(N__17462),
            .I(\Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2 ));
    LocalMux I__4080 (
            .O(N__17459),
            .I(\Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2 ));
    InMux I__4079 (
            .O(N__17454),
            .I(N__17446));
    InMux I__4078 (
            .O(N__17453),
            .I(N__17443));
    InMux I__4077 (
            .O(N__17452),
            .I(N__17436));
    InMux I__4076 (
            .O(N__17451),
            .I(N__17436));
    InMux I__4075 (
            .O(N__17450),
            .I(N__17436));
    InMux I__4074 (
            .O(N__17449),
            .I(N__17433));
    LocalMux I__4073 (
            .O(N__17446),
            .I(N__17430));
    LocalMux I__4072 (
            .O(N__17443),
            .I(N__17425));
    LocalMux I__4071 (
            .O(N__17436),
            .I(N__17425));
    LocalMux I__4070 (
            .O(N__17433),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    Odrv12 I__4069 (
            .O(N__17430),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    Odrv4 I__4068 (
            .O(N__17425),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    CascadeMux I__4067 (
            .O(N__17418),
            .I(\buart.Z_rx.valid_0_cascade_ ));
    CascadeMux I__4066 (
            .O(N__17415),
            .I(N__17412));
    InMux I__4065 (
            .O(N__17412),
            .I(N__17406));
    InMux I__4064 (
            .O(N__17411),
            .I(N__17399));
    InMux I__4063 (
            .O(N__17410),
            .I(N__17399));
    InMux I__4062 (
            .O(N__17409),
            .I(N__17396));
    LocalMux I__4061 (
            .O(N__17406),
            .I(N__17393));
    InMux I__4060 (
            .O(N__17405),
            .I(N__17390));
    InMux I__4059 (
            .O(N__17404),
            .I(N__17387));
    LocalMux I__4058 (
            .O(N__17399),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__4057 (
            .O(N__17396),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    Odrv4 I__4056 (
            .O(N__17393),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__4055 (
            .O(N__17390),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__4054 (
            .O(N__17387),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    CascadeMux I__4053 (
            .O(N__17376),
            .I(bu_rx_data_rdy_cascade_));
    CascadeMux I__4052 (
            .O(N__17373),
            .I(N__17369));
    InMux I__4051 (
            .O(N__17372),
            .I(N__17361));
    InMux I__4050 (
            .O(N__17369),
            .I(N__17361));
    InMux I__4049 (
            .O(N__17368),
            .I(N__17358));
    InMux I__4048 (
            .O(N__17367),
            .I(N__17353));
    InMux I__4047 (
            .O(N__17366),
            .I(N__17353));
    LocalMux I__4046 (
            .O(N__17361),
            .I(N__17350));
    LocalMux I__4045 (
            .O(N__17358),
            .I(N__17345));
    LocalMux I__4044 (
            .O(N__17353),
            .I(N__17345));
    Odrv12 I__4043 (
            .O(N__17350),
            .I(\buart.Z_rx.N_27_0_i ));
    Odrv4 I__4042 (
            .O(N__17345),
            .I(\buart.Z_rx.N_27_0_i ));
    InMux I__4041 (
            .O(N__17340),
            .I(N__17334));
    InMux I__4040 (
            .O(N__17339),
            .I(N__17331));
    InMux I__4039 (
            .O(N__17338),
            .I(N__17326));
    InMux I__4038 (
            .O(N__17337),
            .I(N__17326));
    LocalMux I__4037 (
            .O(N__17334),
            .I(N__17323));
    LocalMux I__4036 (
            .O(N__17331),
            .I(N__17318));
    LocalMux I__4035 (
            .O(N__17326),
            .I(N__17318));
    Odrv12 I__4034 (
            .O(N__17323),
            .I(\Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1 ));
    Odrv4 I__4033 (
            .O(N__17318),
            .I(\Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1 ));
    InMux I__4032 (
            .O(N__17313),
            .I(N__17310));
    LocalMux I__4031 (
            .O(N__17310),
            .I(\Lab_UT.dictrl.next_state_out_2 ));
    InMux I__4030 (
            .O(N__17307),
            .I(N__17302));
    CascadeMux I__4029 (
            .O(N__17306),
            .I(N__17299));
    CascadeMux I__4028 (
            .O(N__17305),
            .I(N__17295));
    LocalMux I__4027 (
            .O(N__17302),
            .I(N__17292));
    InMux I__4026 (
            .O(N__17299),
            .I(N__17289));
    InMux I__4025 (
            .O(N__17298),
            .I(N__17286));
    InMux I__4024 (
            .O(N__17295),
            .I(N__17283));
    Odrv4 I__4023 (
            .O(N__17292),
            .I(\Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ));
    LocalMux I__4022 (
            .O(N__17289),
            .I(\Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ));
    LocalMux I__4021 (
            .O(N__17286),
            .I(\Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ));
    LocalMux I__4020 (
            .O(N__17283),
            .I(\Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ));
    CascadeMux I__4019 (
            .O(N__17274),
            .I(N__17270));
    CascadeMux I__4018 (
            .O(N__17273),
            .I(N__17264));
    InMux I__4017 (
            .O(N__17270),
            .I(N__17261));
    InMux I__4016 (
            .O(N__17269),
            .I(N__17258));
    InMux I__4015 (
            .O(N__17268),
            .I(N__17253));
    InMux I__4014 (
            .O(N__17267),
            .I(N__17253));
    InMux I__4013 (
            .O(N__17264),
            .I(N__17250));
    LocalMux I__4012 (
            .O(N__17261),
            .I(N__17247));
    LocalMux I__4011 (
            .O(N__17258),
            .I(N__17242));
    LocalMux I__4010 (
            .O(N__17253),
            .I(N__17242));
    LocalMux I__4009 (
            .O(N__17250),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    Odrv4 I__4008 (
            .O(N__17247),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    Odrv12 I__4007 (
            .O(N__17242),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__4006 (
            .O(N__17235),
            .I(N__17231));
    InMux I__4005 (
            .O(N__17234),
            .I(N__17224));
    InMux I__4004 (
            .O(N__17231),
            .I(N__17219));
    InMux I__4003 (
            .O(N__17230),
            .I(N__17219));
    InMux I__4002 (
            .O(N__17229),
            .I(N__17214));
    InMux I__4001 (
            .O(N__17228),
            .I(N__17214));
    InMux I__4000 (
            .O(N__17227),
            .I(N__17211));
    LocalMux I__3999 (
            .O(N__17224),
            .I(N__17204));
    LocalMux I__3998 (
            .O(N__17219),
            .I(N__17204));
    LocalMux I__3997 (
            .O(N__17214),
            .I(N__17204));
    LocalMux I__3996 (
            .O(N__17211),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv12 I__3995 (
            .O(N__17204),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    CascadeMux I__3994 (
            .O(N__17199),
            .I(N__17193));
    CascadeMux I__3993 (
            .O(N__17198),
            .I(N__17190));
    CascadeMux I__3992 (
            .O(N__17197),
            .I(N__17187));
    CascadeMux I__3991 (
            .O(N__17196),
            .I(N__17183));
    InMux I__3990 (
            .O(N__17193),
            .I(N__17179));
    InMux I__3989 (
            .O(N__17190),
            .I(N__17176));
    InMux I__3988 (
            .O(N__17187),
            .I(N__17173));
    InMux I__3987 (
            .O(N__17186),
            .I(N__17168));
    InMux I__3986 (
            .O(N__17183),
            .I(N__17168));
    CascadeMux I__3985 (
            .O(N__17182),
            .I(N__17165));
    LocalMux I__3984 (
            .O(N__17179),
            .I(N__17156));
    LocalMux I__3983 (
            .O(N__17176),
            .I(N__17156));
    LocalMux I__3982 (
            .O(N__17173),
            .I(N__17156));
    LocalMux I__3981 (
            .O(N__17168),
            .I(N__17156));
    InMux I__3980 (
            .O(N__17165),
            .I(N__17153));
    Span4Mux_v I__3979 (
            .O(N__17156),
            .I(N__17150));
    LocalMux I__3978 (
            .O(N__17153),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    Odrv4 I__3977 (
            .O(N__17150),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    InMux I__3976 (
            .O(N__17145),
            .I(N__17142));
    LocalMux I__3975 (
            .O(N__17142),
            .I(\buart.Z_rx.idle_0 ));
    InMux I__3974 (
            .O(N__17139),
            .I(N__17135));
    InMux I__3973 (
            .O(N__17138),
            .I(N__17132));
    LocalMux I__3972 (
            .O(N__17135),
            .I(\buart.Z_rx.idle ));
    LocalMux I__3971 (
            .O(N__17132),
            .I(\buart.Z_rx.idle ));
    InMux I__3970 (
            .O(N__17127),
            .I(N__17124));
    LocalMux I__3969 (
            .O(N__17124),
            .I(N__17118));
    InMux I__3968 (
            .O(N__17123),
            .I(N__17115));
    InMux I__3967 (
            .O(N__17122),
            .I(N__17110));
    InMux I__3966 (
            .O(N__17121),
            .I(N__17110));
    Span4Mux_v I__3965 (
            .O(N__17118),
            .I(N__17105));
    LocalMux I__3964 (
            .O(N__17115),
            .I(N__17105));
    LocalMux I__3963 (
            .O(N__17110),
            .I(\buart.Z_rx.ser_clk_2 ));
    Odrv4 I__3962 (
            .O(N__17105),
            .I(\buart.Z_rx.ser_clk_2 ));
    CascadeMux I__3961 (
            .O(N__17100),
            .I(N__17095));
    InMux I__3960 (
            .O(N__17099),
            .I(N__17091));
    InMux I__3959 (
            .O(N__17098),
            .I(N__17088));
    InMux I__3958 (
            .O(N__17095),
            .I(N__17084));
    InMux I__3957 (
            .O(N__17094),
            .I(N__17081));
    LocalMux I__3956 (
            .O(N__17091),
            .I(N__17076));
    LocalMux I__3955 (
            .O(N__17088),
            .I(N__17076));
    InMux I__3954 (
            .O(N__17087),
            .I(N__17073));
    LocalMux I__3953 (
            .O(N__17084),
            .I(N__17066));
    LocalMux I__3952 (
            .O(N__17081),
            .I(N__17066));
    Span4Mux_v I__3951 (
            .O(N__17076),
            .I(N__17066));
    LocalMux I__3950 (
            .O(N__17073),
            .I(\buart.Z_rx.ser_clk_3 ));
    Odrv4 I__3949 (
            .O(N__17066),
            .I(\buart.Z_rx.ser_clk_3 ));
    CascadeMux I__3948 (
            .O(N__17061),
            .I(\buart.Z_rx.idle_cascade_ ));
    InMux I__3947 (
            .O(N__17058),
            .I(N__17055));
    LocalMux I__3946 (
            .O(N__17055),
            .I(N__17051));
    InMux I__3945 (
            .O(N__17054),
            .I(N__17048));
    Span4Mux_h I__3944 (
            .O(N__17051),
            .I(N__17045));
    LocalMux I__3943 (
            .O(N__17048),
            .I(bu_rx_data_rdy));
    Odrv4 I__3942 (
            .O(N__17045),
            .I(bu_rx_data_rdy));
    CascadeMux I__3941 (
            .O(N__17040),
            .I(N__17034));
    CascadeMux I__3940 (
            .O(N__17039),
            .I(N__17031));
    InMux I__3939 (
            .O(N__17038),
            .I(N__17022));
    InMux I__3938 (
            .O(N__17037),
            .I(N__17022));
    InMux I__3937 (
            .O(N__17034),
            .I(N__17022));
    InMux I__3936 (
            .O(N__17031),
            .I(N__17022));
    LocalMux I__3935 (
            .O(N__17022),
            .I(N__17018));
    InMux I__3934 (
            .O(N__17021),
            .I(N__17015));
    Odrv12 I__3933 (
            .O(N__17018),
            .I(\buart.Z_rx.bitcountlde_0 ));
    LocalMux I__3932 (
            .O(N__17015),
            .I(\buart.Z_rx.bitcountlde_0 ));
    InMux I__3931 (
            .O(N__17010),
            .I(N__17007));
    LocalMux I__3930 (
            .O(N__17007),
            .I(N__17003));
    InMux I__3929 (
            .O(N__17006),
            .I(N__16999));
    Span4Mux_h I__3928 (
            .O(N__17003),
            .I(N__16995));
    InMux I__3927 (
            .O(N__17002),
            .I(N__16992));
    LocalMux I__3926 (
            .O(N__16999),
            .I(N__16989));
    InMux I__3925 (
            .O(N__16998),
            .I(N__16986));
    Odrv4 I__3924 (
            .O(N__16995),
            .I(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ));
    LocalMux I__3923 (
            .O(N__16992),
            .I(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ));
    Odrv4 I__3922 (
            .O(N__16989),
            .I(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ));
    LocalMux I__3921 (
            .O(N__16986),
            .I(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ));
    CascadeMux I__3920 (
            .O(N__16977),
            .I(N__16973));
    InMux I__3919 (
            .O(N__16976),
            .I(N__16969));
    InMux I__3918 (
            .O(N__16973),
            .I(N__16966));
    InMux I__3917 (
            .O(N__16972),
            .I(N__16963));
    LocalMux I__3916 (
            .O(N__16969),
            .I(N__16960));
    LocalMux I__3915 (
            .O(N__16966),
            .I(N__16956));
    LocalMux I__3914 (
            .O(N__16963),
            .I(N__16953));
    Span4Mux_h I__3913 (
            .O(N__16960),
            .I(N__16950));
    InMux I__3912 (
            .O(N__16959),
            .I(N__16947));
    Odrv4 I__3911 (
            .O(N__16956),
            .I(\Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ));
    Odrv4 I__3910 (
            .O(N__16953),
            .I(\Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ));
    Odrv4 I__3909 (
            .O(N__16950),
            .I(\Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ));
    LocalMux I__3908 (
            .O(N__16947),
            .I(\Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ));
    InMux I__3907 (
            .O(N__16938),
            .I(N__16932));
    InMux I__3906 (
            .O(N__16937),
            .I(N__16929));
    InMux I__3905 (
            .O(N__16936),
            .I(N__16926));
    InMux I__3904 (
            .O(N__16935),
            .I(N__16923));
    LocalMux I__3903 (
            .O(N__16932),
            .I(N__16920));
    LocalMux I__3902 (
            .O(N__16929),
            .I(N__16915));
    LocalMux I__3901 (
            .O(N__16926),
            .I(N__16915));
    LocalMux I__3900 (
            .O(N__16923),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    Odrv4 I__3899 (
            .O(N__16920),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    Odrv4 I__3898 (
            .O(N__16915),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    InMux I__3897 (
            .O(N__16908),
            .I(N__16900));
    InMux I__3896 (
            .O(N__16907),
            .I(N__16900));
    InMux I__3895 (
            .O(N__16906),
            .I(N__16897));
    InMux I__3894 (
            .O(N__16905),
            .I(N__16894));
    LocalMux I__3893 (
            .O(N__16900),
            .I(N__16890));
    LocalMux I__3892 (
            .O(N__16897),
            .I(N__16885));
    LocalMux I__3891 (
            .O(N__16894),
            .I(N__16885));
    CascadeMux I__3890 (
            .O(N__16893),
            .I(N__16879));
    Span4Mux_h I__3889 (
            .O(N__16890),
            .I(N__16874));
    Span4Mux_s3_v I__3888 (
            .O(N__16885),
            .I(N__16871));
    InMux I__3887 (
            .O(N__16884),
            .I(N__16864));
    InMux I__3886 (
            .O(N__16883),
            .I(N__16864));
    InMux I__3885 (
            .O(N__16882),
            .I(N__16864));
    InMux I__3884 (
            .O(N__16879),
            .I(N__16857));
    InMux I__3883 (
            .O(N__16878),
            .I(N__16857));
    InMux I__3882 (
            .O(N__16877),
            .I(N__16857));
    Odrv4 I__3881 (
            .O(N__16874),
            .I(\Lab_UT.state_i_3_3 ));
    Odrv4 I__3880 (
            .O(N__16871),
            .I(\Lab_UT.state_i_3_3 ));
    LocalMux I__3879 (
            .O(N__16864),
            .I(\Lab_UT.state_i_3_3 ));
    LocalMux I__3878 (
            .O(N__16857),
            .I(\Lab_UT.state_i_3_3 ));
    InMux I__3877 (
            .O(N__16848),
            .I(N__16845));
    LocalMux I__3876 (
            .O(N__16845),
            .I(N__16841));
    InMux I__3875 (
            .O(N__16844),
            .I(N__16838));
    Odrv4 I__3874 (
            .O(N__16841),
            .I(\Lab_UT.alarmcharZ0Z_1 ));
    LocalMux I__3873 (
            .O(N__16838),
            .I(\Lab_UT.alarmcharZ0Z_1 ));
    InMux I__3872 (
            .O(N__16833),
            .I(N__16829));
    InMux I__3871 (
            .O(N__16832),
            .I(N__16818));
    LocalMux I__3870 (
            .O(N__16829),
            .I(N__16813));
    CascadeMux I__3869 (
            .O(N__16828),
            .I(N__16807));
    InMux I__3868 (
            .O(N__16827),
            .I(N__16800));
    InMux I__3867 (
            .O(N__16826),
            .I(N__16800));
    InMux I__3866 (
            .O(N__16825),
            .I(N__16800));
    InMux I__3865 (
            .O(N__16824),
            .I(N__16795));
    InMux I__3864 (
            .O(N__16823),
            .I(N__16795));
    CascadeMux I__3863 (
            .O(N__16822),
            .I(N__16791));
    InMux I__3862 (
            .O(N__16821),
            .I(N__16787));
    LocalMux I__3861 (
            .O(N__16818),
            .I(N__16784));
    InMux I__3860 (
            .O(N__16817),
            .I(N__16779));
    InMux I__3859 (
            .O(N__16816),
            .I(N__16779));
    Span4Mux_v I__3858 (
            .O(N__16813),
            .I(N__16776));
    InMux I__3857 (
            .O(N__16812),
            .I(N__16773));
    InMux I__3856 (
            .O(N__16811),
            .I(N__16768));
    InMux I__3855 (
            .O(N__16810),
            .I(N__16768));
    InMux I__3854 (
            .O(N__16807),
            .I(N__16765));
    LocalMux I__3853 (
            .O(N__16800),
            .I(N__16760));
    LocalMux I__3852 (
            .O(N__16795),
            .I(N__16760));
    InMux I__3851 (
            .O(N__16794),
            .I(N__16753));
    InMux I__3850 (
            .O(N__16791),
            .I(N__16753));
    InMux I__3849 (
            .O(N__16790),
            .I(N__16753));
    LocalMux I__3848 (
            .O(N__16787),
            .I(N__16750));
    Span4Mux_h I__3847 (
            .O(N__16784),
            .I(N__16747));
    LocalMux I__3846 (
            .O(N__16779),
            .I(\Lab_UT.cnt_3 ));
    Odrv4 I__3845 (
            .O(N__16776),
            .I(\Lab_UT.cnt_3 ));
    LocalMux I__3844 (
            .O(N__16773),
            .I(\Lab_UT.cnt_3 ));
    LocalMux I__3843 (
            .O(N__16768),
            .I(\Lab_UT.cnt_3 ));
    LocalMux I__3842 (
            .O(N__16765),
            .I(\Lab_UT.cnt_3 ));
    Odrv4 I__3841 (
            .O(N__16760),
            .I(\Lab_UT.cnt_3 ));
    LocalMux I__3840 (
            .O(N__16753),
            .I(\Lab_UT.cnt_3 ));
    Odrv12 I__3839 (
            .O(N__16750),
            .I(\Lab_UT.cnt_3 ));
    Odrv4 I__3838 (
            .O(N__16747),
            .I(\Lab_UT.cnt_3 ));
    CascadeMux I__3837 (
            .O(N__16728),
            .I(N__16725));
    InMux I__3836 (
            .O(N__16725),
            .I(N__16715));
    CascadeMux I__3835 (
            .O(N__16724),
            .I(N__16712));
    InMux I__3834 (
            .O(N__16723),
            .I(N__16707));
    CascadeMux I__3833 (
            .O(N__16722),
            .I(N__16702));
    CascadeMux I__3832 (
            .O(N__16721),
            .I(N__16699));
    CascadeMux I__3831 (
            .O(N__16720),
            .I(N__16696));
    InMux I__3830 (
            .O(N__16719),
            .I(N__16689));
    InMux I__3829 (
            .O(N__16718),
            .I(N__16689));
    LocalMux I__3828 (
            .O(N__16715),
            .I(N__16686));
    InMux I__3827 (
            .O(N__16712),
            .I(N__16678));
    InMux I__3826 (
            .O(N__16711),
            .I(N__16678));
    InMux I__3825 (
            .O(N__16710),
            .I(N__16678));
    LocalMux I__3824 (
            .O(N__16707),
            .I(N__16675));
    InMux I__3823 (
            .O(N__16706),
            .I(N__16668));
    InMux I__3822 (
            .O(N__16705),
            .I(N__16668));
    InMux I__3821 (
            .O(N__16702),
            .I(N__16668));
    InMux I__3820 (
            .O(N__16699),
            .I(N__16661));
    InMux I__3819 (
            .O(N__16696),
            .I(N__16661));
    InMux I__3818 (
            .O(N__16695),
            .I(N__16661));
    InMux I__3817 (
            .O(N__16694),
            .I(N__16658));
    LocalMux I__3816 (
            .O(N__16689),
            .I(N__16655));
    Span4Mux_v I__3815 (
            .O(N__16686),
            .I(N__16652));
    InMux I__3814 (
            .O(N__16685),
            .I(N__16649));
    LocalMux I__3813 (
            .O(N__16678),
            .I(N__16640));
    Sp12to4 I__3812 (
            .O(N__16675),
            .I(N__16640));
    LocalMux I__3811 (
            .O(N__16668),
            .I(N__16640));
    LocalMux I__3810 (
            .O(N__16661),
            .I(N__16640));
    LocalMux I__3809 (
            .O(N__16658),
            .I(N__16633));
    Span4Mux_v I__3808 (
            .O(N__16655),
            .I(N__16633));
    Span4Mux_h I__3807 (
            .O(N__16652),
            .I(N__16633));
    LocalMux I__3806 (
            .O(N__16649),
            .I(\Lab_UT.cnt_1 ));
    Odrv12 I__3805 (
            .O(N__16640),
            .I(\Lab_UT.cnt_1 ));
    Odrv4 I__3804 (
            .O(N__16633),
            .I(\Lab_UT.cnt_1 ));
    InMux I__3803 (
            .O(N__16626),
            .I(N__16623));
    LocalMux I__3802 (
            .O(N__16623),
            .I(N__16620));
    Span4Mux_h I__3801 (
            .O(N__16620),
            .I(N__16617));
    Odrv4 I__3800 (
            .O(N__16617),
            .I(\Lab_UT.bcd2segment1.m42_bmZ0 ));
    IoInMux I__3799 (
            .O(N__16614),
            .I(N__16611));
    LocalMux I__3798 (
            .O(N__16611),
            .I(N__16608));
    IoSpan4Mux I__3797 (
            .O(N__16608),
            .I(N__16603));
    SRMux I__3796 (
            .O(N__16607),
            .I(N__16600));
    InMux I__3795 (
            .O(N__16606),
            .I(N__16596));
    Span4Mux_s1_v I__3794 (
            .O(N__16603),
            .I(N__16593));
    LocalMux I__3793 (
            .O(N__16600),
            .I(N__16590));
    InMux I__3792 (
            .O(N__16599),
            .I(N__16587));
    LocalMux I__3791 (
            .O(N__16596),
            .I(N__16584));
    Span4Mux_v I__3790 (
            .O(N__16593),
            .I(N__16579));
    Span4Mux_s3_h I__3789 (
            .O(N__16590),
            .I(N__16579));
    LocalMux I__3788 (
            .O(N__16587),
            .I(N__16576));
    Span12Mux_s6_h I__3787 (
            .O(N__16584),
            .I(N__16573));
    Span4Mux_h I__3786 (
            .O(N__16579),
            .I(N__16568));
    Span4Mux_h I__3785 (
            .O(N__16576),
            .I(N__16568));
    Odrv12 I__3784 (
            .O(N__16573),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3783 (
            .O(N__16568),
            .I(CONSTANT_ONE_NET));
    InMux I__3782 (
            .O(N__16563),
            .I(N__16560));
    LocalMux I__3781 (
            .O(N__16560),
            .I(N__16557));
    Odrv4 I__3780 (
            .O(N__16557),
            .I(\buart.Z_rx.bitcount_lm_0 ));
    CascadeMux I__3779 (
            .O(N__16554),
            .I(\buart.Z_rx.un1_sample_0_cascade_ ));
    InMux I__3778 (
            .O(N__16551),
            .I(N__16548));
    LocalMux I__3777 (
            .O(N__16548),
            .I(N__16545));
    Odrv4 I__3776 (
            .O(N__16545),
            .I(\Lab_UT.dictrl.next_state_out_3 ));
    SRMux I__3775 (
            .O(N__16542),
            .I(N__16539));
    LocalMux I__3774 (
            .O(N__16539),
            .I(N__16536));
    Span4Mux_h I__3773 (
            .O(N__16536),
            .I(N__16533));
    Odrv4 I__3772 (
            .O(N__16533),
            .I(\Lab_UT.m68_0_ns ));
    InMux I__3771 (
            .O(N__16530),
            .I(N__16527));
    LocalMux I__3770 (
            .O(N__16527),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__3769 (
            .O(N__16524),
            .I(N__16521));
    LocalMux I__3768 (
            .O(N__16521),
            .I(N__16518));
    Odrv12 I__3767 (
            .O(N__16518),
            .I(\buart.Z_rx.bitcount_lm_1 ));
    InMux I__3766 (
            .O(N__16515),
            .I(N__16506));
    InMux I__3765 (
            .O(N__16514),
            .I(N__16501));
    InMux I__3764 (
            .O(N__16513),
            .I(N__16501));
    InMux I__3763 (
            .O(N__16512),
            .I(N__16492));
    InMux I__3762 (
            .O(N__16511),
            .I(N__16492));
    InMux I__3761 (
            .O(N__16510),
            .I(N__16492));
    InMux I__3760 (
            .O(N__16509),
            .I(N__16492));
    LocalMux I__3759 (
            .O(N__16506),
            .I(N__16480));
    LocalMux I__3758 (
            .O(N__16501),
            .I(N__16477));
    LocalMux I__3757 (
            .O(N__16492),
            .I(N__16474));
    InMux I__3756 (
            .O(N__16491),
            .I(N__16469));
    InMux I__3755 (
            .O(N__16490),
            .I(N__16469));
    InMux I__3754 (
            .O(N__16489),
            .I(N__16464));
    InMux I__3753 (
            .O(N__16488),
            .I(N__16464));
    InMux I__3752 (
            .O(N__16487),
            .I(N__16461));
    InMux I__3751 (
            .O(N__16486),
            .I(N__16456));
    InMux I__3750 (
            .O(N__16485),
            .I(N__16456));
    InMux I__3749 (
            .O(N__16484),
            .I(N__16451));
    InMux I__3748 (
            .O(N__16483),
            .I(N__16451));
    Span4Mux_h I__3747 (
            .O(N__16480),
            .I(N__16448));
    Span4Mux_h I__3746 (
            .O(N__16477),
            .I(N__16443));
    Span4Mux_v I__3745 (
            .O(N__16474),
            .I(N__16443));
    LocalMux I__3744 (
            .O(N__16469),
            .I(N__16438));
    LocalMux I__3743 (
            .O(N__16464),
            .I(N__16438));
    LocalMux I__3742 (
            .O(N__16461),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__3741 (
            .O(N__16456),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__3740 (
            .O(N__16451),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__3739 (
            .O(N__16448),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__3738 (
            .O(N__16443),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__3737 (
            .O(N__16438),
            .I(\buart.Z_rx.startbit ));
    InMux I__3736 (
            .O(N__16425),
            .I(N__16422));
    LocalMux I__3735 (
            .O(N__16422),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__3734 (
            .O(N__16419),
            .I(N__16416));
    LocalMux I__3733 (
            .O(N__16416),
            .I(N__16413));
    Odrv12 I__3732 (
            .O(N__16413),
            .I(\buart.Z_rx.bitcount_lm_2 ));
    CascadeMux I__3731 (
            .O(N__16410),
            .I(N__16405));
    CascadeMux I__3730 (
            .O(N__16409),
            .I(N__16402));
    CascadeMux I__3729 (
            .O(N__16408),
            .I(N__16399));
    InMux I__3728 (
            .O(N__16405),
            .I(N__16388));
    InMux I__3727 (
            .O(N__16402),
            .I(N__16388));
    InMux I__3726 (
            .O(N__16399),
            .I(N__16388));
    InMux I__3725 (
            .O(N__16398),
            .I(N__16388));
    InMux I__3724 (
            .O(N__16397),
            .I(N__16384));
    LocalMux I__3723 (
            .O(N__16388),
            .I(N__16379));
    CascadeMux I__3722 (
            .O(N__16387),
            .I(N__16375));
    LocalMux I__3721 (
            .O(N__16384),
            .I(N__16370));
    CascadeMux I__3720 (
            .O(N__16383),
            .I(N__16367));
    CascadeMux I__3719 (
            .O(N__16382),
            .I(N__16364));
    Span4Mux_s2_v I__3718 (
            .O(N__16379),
            .I(N__16357));
    InMux I__3717 (
            .O(N__16378),
            .I(N__16354));
    InMux I__3716 (
            .O(N__16375),
            .I(N__16351));
    InMux I__3715 (
            .O(N__16374),
            .I(N__16346));
    InMux I__3714 (
            .O(N__16373),
            .I(N__16346));
    Span4Mux_h I__3713 (
            .O(N__16370),
            .I(N__16343));
    InMux I__3712 (
            .O(N__16367),
            .I(N__16336));
    InMux I__3711 (
            .O(N__16364),
            .I(N__16336));
    InMux I__3710 (
            .O(N__16363),
            .I(N__16336));
    InMux I__3709 (
            .O(N__16362),
            .I(N__16329));
    InMux I__3708 (
            .O(N__16361),
            .I(N__16329));
    InMux I__3707 (
            .O(N__16360),
            .I(N__16329));
    Span4Mux_v I__3706 (
            .O(N__16357),
            .I(N__16326));
    LocalMux I__3705 (
            .O(N__16354),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3704 (
            .O(N__16351),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3703 (
            .O(N__16346),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__3702 (
            .O(N__16343),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3701 (
            .O(N__16336),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3700 (
            .O(N__16329),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__3699 (
            .O(N__16326),
            .I(\Lab_UT.di_Mtens_0 ));
    InMux I__3698 (
            .O(N__16311),
            .I(N__16308));
    LocalMux I__3697 (
            .O(N__16308),
            .I(N__16305));
    Odrv12 I__3696 (
            .O(N__16305),
            .I(\Lab_UT.bcd2segment1.N_166 ));
    InMux I__3695 (
            .O(N__16302),
            .I(N__16299));
    LocalMux I__3694 (
            .O(N__16299),
            .I(N__16296));
    Span4Mux_h I__3693 (
            .O(N__16296),
            .I(N__16292));
    CascadeMux I__3692 (
            .O(N__16295),
            .I(N__16289));
    Span4Mux_v I__3691 (
            .O(N__16292),
            .I(N__16285));
    InMux I__3690 (
            .O(N__16289),
            .I(N__16280));
    InMux I__3689 (
            .O(N__16288),
            .I(N__16280));
    Span4Mux_s2_h I__3688 (
            .O(N__16285),
            .I(N__16276));
    LocalMux I__3687 (
            .O(N__16280),
            .I(N__16273));
    InMux I__3686 (
            .O(N__16279),
            .I(N__16270));
    Odrv4 I__3685 (
            .O(N__16276),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    Odrv4 I__3684 (
            .O(N__16273),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    LocalMux I__3683 (
            .O(N__16270),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__3682 (
            .O(N__16263),
            .I(N__16257));
    InMux I__3681 (
            .O(N__16262),
            .I(N__16257));
    LocalMux I__3680 (
            .O(N__16257),
            .I(N__16249));
    InMux I__3679 (
            .O(N__16256),
            .I(N__16244));
    InMux I__3678 (
            .O(N__16255),
            .I(N__16244));
    InMux I__3677 (
            .O(N__16254),
            .I(N__16238));
    InMux I__3676 (
            .O(N__16253),
            .I(N__16235));
    InMux I__3675 (
            .O(N__16252),
            .I(N__16232));
    Span4Mux_h I__3674 (
            .O(N__16249),
            .I(N__16226));
    LocalMux I__3673 (
            .O(N__16244),
            .I(N__16223));
    InMux I__3672 (
            .O(N__16243),
            .I(N__16218));
    InMux I__3671 (
            .O(N__16242),
            .I(N__16218));
    InMux I__3670 (
            .O(N__16241),
            .I(N__16215));
    LocalMux I__3669 (
            .O(N__16238),
            .I(N__16209));
    LocalMux I__3668 (
            .O(N__16235),
            .I(N__16209));
    LocalMux I__3667 (
            .O(N__16232),
            .I(N__16206));
    InMux I__3666 (
            .O(N__16231),
            .I(N__16199));
    InMux I__3665 (
            .O(N__16230),
            .I(N__16199));
    InMux I__3664 (
            .O(N__16229),
            .I(N__16199));
    Span4Mux_v I__3663 (
            .O(N__16226),
            .I(N__16196));
    Span4Mux_v I__3662 (
            .O(N__16223),
            .I(N__16193));
    LocalMux I__3661 (
            .O(N__16218),
            .I(N__16190));
    LocalMux I__3660 (
            .O(N__16215),
            .I(N__16187));
    InMux I__3659 (
            .O(N__16214),
            .I(N__16184));
    Odrv4 I__3658 (
            .O(N__16209),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3657 (
            .O(N__16206),
            .I(\Lab_UT.di_Mones_2 ));
    LocalMux I__3656 (
            .O(N__16199),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3655 (
            .O(N__16196),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3654 (
            .O(N__16193),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3653 (
            .O(N__16190),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv12 I__3652 (
            .O(N__16187),
            .I(\Lab_UT.di_Mones_2 ));
    LocalMux I__3651 (
            .O(N__16184),
            .I(\Lab_UT.di_Mones_2 ));
    InMux I__3650 (
            .O(N__16167),
            .I(N__16164));
    LocalMux I__3649 (
            .O(N__16164),
            .I(N__16161));
    Span4Mux_h I__3648 (
            .O(N__16161),
            .I(N__16158));
    Odrv4 I__3647 (
            .O(N__16158),
            .I(\Lab_UT.didp.countrce3.q_RNO_0Z0Z_3 ));
    InMux I__3646 (
            .O(N__16155),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__3645 (
            .O(N__16152),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    CascadeMux I__3644 (
            .O(N__16149),
            .I(N__16146));
    InMux I__3643 (
            .O(N__16146),
            .I(N__16143));
    LocalMux I__3642 (
            .O(N__16143),
            .I(N__16140));
    Span4Mux_v I__3641 (
            .O(N__16140),
            .I(N__16137));
    Odrv4 I__3640 (
            .O(N__16137),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__3639 (
            .O(N__16134),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__3638 (
            .O(N__16131),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    InMux I__3637 (
            .O(N__16128),
            .I(N__16125));
    LocalMux I__3636 (
            .O(N__16125),
            .I(N__16122));
    Odrv4 I__3635 (
            .O(N__16122),
            .I(\buart.Z_rx.bitcount_lm_4 ));
    InMux I__3634 (
            .O(N__16119),
            .I(N__16112));
    InMux I__3633 (
            .O(N__16118),
            .I(N__16109));
    CascadeMux I__3632 (
            .O(N__16117),
            .I(N__16105));
    CascadeMux I__3631 (
            .O(N__16116),
            .I(N__16099));
    InMux I__3630 (
            .O(N__16115),
            .I(N__16096));
    LocalMux I__3629 (
            .O(N__16112),
            .I(N__16093));
    LocalMux I__3628 (
            .O(N__16109),
            .I(N__16090));
    InMux I__3627 (
            .O(N__16108),
            .I(N__16087));
    InMux I__3626 (
            .O(N__16105),
            .I(N__16080));
    InMux I__3625 (
            .O(N__16104),
            .I(N__16080));
    InMux I__3624 (
            .O(N__16103),
            .I(N__16080));
    InMux I__3623 (
            .O(N__16102),
            .I(N__16077));
    InMux I__3622 (
            .O(N__16099),
            .I(N__16074));
    LocalMux I__3621 (
            .O(N__16096),
            .I(N__16069));
    Span4Mux_h I__3620 (
            .O(N__16093),
            .I(N__16069));
    Span4Mux_h I__3619 (
            .O(N__16090),
            .I(N__16064));
    LocalMux I__3618 (
            .O(N__16087),
            .I(N__16064));
    LocalMux I__3617 (
            .O(N__16080),
            .I(N__16059));
    LocalMux I__3616 (
            .O(N__16077),
            .I(N__16059));
    LocalMux I__3615 (
            .O(N__16074),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    Odrv4 I__3614 (
            .O(N__16069),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    Odrv4 I__3613 (
            .O(N__16064),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    Odrv4 I__3612 (
            .O(N__16059),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    CascadeMux I__3611 (
            .O(N__16050),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_ ));
    InMux I__3610 (
            .O(N__16047),
            .I(N__16044));
    LocalMux I__3609 (
            .O(N__16044),
            .I(\uu2.mem0.N_294 ));
    InMux I__3608 (
            .O(N__16041),
            .I(N__16038));
    LocalMux I__3607 (
            .O(N__16038),
            .I(N__16034));
    InMux I__3606 (
            .O(N__16037),
            .I(N__16031));
    Odrv4 I__3605 (
            .O(N__16034),
            .I(\uu2.bitmapZ0Z_180 ));
    LocalMux I__3604 (
            .O(N__16031),
            .I(\uu2.bitmapZ0Z_180 ));
    InMux I__3603 (
            .O(N__16026),
            .I(N__16023));
    LocalMux I__3602 (
            .O(N__16023),
            .I(\uu2.mem0.N_271 ));
    InMux I__3601 (
            .O(N__16020),
            .I(N__16017));
    LocalMux I__3600 (
            .O(N__16017),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_80 ));
    InMux I__3599 (
            .O(N__16014),
            .I(N__16011));
    LocalMux I__3598 (
            .O(N__16011),
            .I(N__16008));
    Span4Mux_h I__3597 (
            .O(N__16008),
            .I(N__16004));
    InMux I__3596 (
            .O(N__16007),
            .I(N__16001));
    Odrv4 I__3595 (
            .O(N__16004),
            .I(\uu2.bitmapZ0Z_197 ));
    LocalMux I__3594 (
            .O(N__16001),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__3593 (
            .O(N__15996),
            .I(N__15987));
    InMux I__3592 (
            .O(N__15995),
            .I(N__15987));
    InMux I__3591 (
            .O(N__15994),
            .I(N__15984));
    CascadeMux I__3590 (
            .O(N__15993),
            .I(N__15978));
    InMux I__3589 (
            .O(N__15992),
            .I(N__15974));
    LocalMux I__3588 (
            .O(N__15987),
            .I(N__15970));
    LocalMux I__3587 (
            .O(N__15984),
            .I(N__15967));
    InMux I__3586 (
            .O(N__15983),
            .I(N__15961));
    InMux I__3585 (
            .O(N__15982),
            .I(N__15961));
    InMux I__3584 (
            .O(N__15981),
            .I(N__15954));
    InMux I__3583 (
            .O(N__15978),
            .I(N__15954));
    InMux I__3582 (
            .O(N__15977),
            .I(N__15954));
    LocalMux I__3581 (
            .O(N__15974),
            .I(N__15951));
    InMux I__3580 (
            .O(N__15973),
            .I(N__15948));
    Span4Mux_v I__3579 (
            .O(N__15970),
            .I(N__15943));
    Span4Mux_v I__3578 (
            .O(N__15967),
            .I(N__15943));
    InMux I__3577 (
            .O(N__15966),
            .I(N__15940));
    LocalMux I__3576 (
            .O(N__15961),
            .I(N__15937));
    LocalMux I__3575 (
            .O(N__15954),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3574 (
            .O(N__15951),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__3573 (
            .O(N__15948),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3572 (
            .O(N__15943),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__3571 (
            .O(N__15940),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3570 (
            .O(N__15937),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    InMux I__3569 (
            .O(N__15924),
            .I(N__15921));
    LocalMux I__3568 (
            .O(N__15921),
            .I(N__15918));
    Span4Mux_v I__3567 (
            .O(N__15918),
            .I(N__15914));
    InMux I__3566 (
            .O(N__15917),
            .I(N__15911));
    Odrv4 I__3565 (
            .O(N__15914),
            .I(\uu2.bitmapZ0Z_69 ));
    LocalMux I__3564 (
            .O(N__15911),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__3563 (
            .O(N__15906),
            .I(N__15903));
    LocalMux I__3562 (
            .O(N__15903),
            .I(N__15900));
    Span4Mux_h I__3561 (
            .O(N__15900),
            .I(N__15897));
    Odrv4 I__3560 (
            .O(N__15897),
            .I(\uu2.mem0.N_98_0 ));
    CascadeMux I__3559 (
            .O(N__15894),
            .I(N__15890));
    InMux I__3558 (
            .O(N__15893),
            .I(N__15886));
    InMux I__3557 (
            .O(N__15890),
            .I(N__15883));
    InMux I__3556 (
            .O(N__15889),
            .I(N__15880));
    LocalMux I__3555 (
            .O(N__15886),
            .I(N__15877));
    LocalMux I__3554 (
            .O(N__15883),
            .I(N__15872));
    LocalMux I__3553 (
            .O(N__15880),
            .I(N__15872));
    Span4Mux_h I__3552 (
            .O(N__15877),
            .I(N__15869));
    Span4Mux_h I__3551 (
            .O(N__15872),
            .I(N__15865));
    Span4Mux_v I__3550 (
            .O(N__15869),
            .I(N__15862));
    InMux I__3549 (
            .O(N__15868),
            .I(N__15859));
    Span4Mux_h I__3548 (
            .O(N__15865),
            .I(N__15856));
    Odrv4 I__3547 (
            .O(N__15862),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__3546 (
            .O(N__15859),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__3545 (
            .O(N__15856),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__3544 (
            .O(N__15849),
            .I(N__15845));
    CascadeMux I__3543 (
            .O(N__15848),
            .I(N__15841));
    InMux I__3542 (
            .O(N__15845),
            .I(N__15836));
    InMux I__3541 (
            .O(N__15844),
            .I(N__15836));
    InMux I__3540 (
            .O(N__15841),
            .I(N__15831));
    LocalMux I__3539 (
            .O(N__15836),
            .I(N__15828));
    InMux I__3538 (
            .O(N__15835),
            .I(N__15825));
    InMux I__3537 (
            .O(N__15834),
            .I(N__15821));
    LocalMux I__3536 (
            .O(N__15831),
            .I(N__15818));
    Span4Mux_h I__3535 (
            .O(N__15828),
            .I(N__15815));
    LocalMux I__3534 (
            .O(N__15825),
            .I(N__15812));
    InMux I__3533 (
            .O(N__15824),
            .I(N__15809));
    LocalMux I__3532 (
            .O(N__15821),
            .I(N__15806));
    Odrv4 I__3531 (
            .O(N__15818),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__3530 (
            .O(N__15815),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv12 I__3529 (
            .O(N__15812),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__3528 (
            .O(N__15809),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__3527 (
            .O(N__15806),
            .I(\uu2.r_addrZ0Z_0 ));
    InMux I__3526 (
            .O(N__15795),
            .I(N__15789));
    InMux I__3525 (
            .O(N__15794),
            .I(N__15789));
    LocalMux I__3524 (
            .O(N__15789),
            .I(N__15782));
    InMux I__3523 (
            .O(N__15788),
            .I(N__15773));
    InMux I__3522 (
            .O(N__15787),
            .I(N__15773));
    InMux I__3521 (
            .O(N__15786),
            .I(N__15773));
    InMux I__3520 (
            .O(N__15785),
            .I(N__15773));
    Odrv12 I__3519 (
            .O(N__15782),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__3518 (
            .O(N__15773),
            .I(\uu2.trig_rd_is_det ));
    InMux I__3517 (
            .O(N__15768),
            .I(N__15765));
    LocalMux I__3516 (
            .O(N__15765),
            .I(N__15761));
    CascadeMux I__3515 (
            .O(N__15764),
            .I(N__15758));
    Span4Mux_v I__3514 (
            .O(N__15761),
            .I(N__15755));
    InMux I__3513 (
            .O(N__15758),
            .I(N__15751));
    IoSpan4Mux I__3512 (
            .O(N__15755),
            .I(N__15748));
    InMux I__3511 (
            .O(N__15754),
            .I(N__15745));
    LocalMux I__3510 (
            .O(N__15751),
            .I(N__15738));
    Span4Mux_s0_h I__3509 (
            .O(N__15748),
            .I(N__15738));
    LocalMux I__3508 (
            .O(N__15745),
            .I(N__15738));
    Span4Mux_h I__3507 (
            .O(N__15738),
            .I(N__15733));
    InMux I__3506 (
            .O(N__15737),
            .I(N__15728));
    InMux I__3505 (
            .O(N__15736),
            .I(N__15728));
    Span4Mux_h I__3504 (
            .O(N__15733),
            .I(N__15725));
    LocalMux I__3503 (
            .O(N__15728),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv4 I__3502 (
            .O(N__15725),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__3501 (
            .O(N__15720),
            .I(\uu2.N_12_i_cascade_ ));
    InMux I__3500 (
            .O(N__15717),
            .I(N__15708));
    InMux I__3499 (
            .O(N__15716),
            .I(N__15701));
    InMux I__3498 (
            .O(N__15715),
            .I(N__15701));
    InMux I__3497 (
            .O(N__15714),
            .I(N__15701));
    InMux I__3496 (
            .O(N__15713),
            .I(N__15698));
    InMux I__3495 (
            .O(N__15712),
            .I(N__15693));
    InMux I__3494 (
            .O(N__15711),
            .I(N__15693));
    LocalMux I__3493 (
            .O(N__15708),
            .I(N__15688));
    LocalMux I__3492 (
            .O(N__15701),
            .I(N__15688));
    LocalMux I__3491 (
            .O(N__15698),
            .I(\uu2.N_67 ));
    LocalMux I__3490 (
            .O(N__15693),
            .I(\uu2.N_67 ));
    Odrv12 I__3489 (
            .O(N__15688),
            .I(\uu2.N_67 ));
    InMux I__3488 (
            .O(N__15681),
            .I(N__15665));
    InMux I__3487 (
            .O(N__15680),
            .I(N__15665));
    InMux I__3486 (
            .O(N__15679),
            .I(N__15665));
    InMux I__3485 (
            .O(N__15678),
            .I(N__15662));
    InMux I__3484 (
            .O(N__15677),
            .I(N__15659));
    InMux I__3483 (
            .O(N__15676),
            .I(N__15654));
    InMux I__3482 (
            .O(N__15675),
            .I(N__15654));
    InMux I__3481 (
            .O(N__15674),
            .I(N__15644));
    InMux I__3480 (
            .O(N__15673),
            .I(N__15644));
    InMux I__3479 (
            .O(N__15672),
            .I(N__15644));
    LocalMux I__3478 (
            .O(N__15665),
            .I(N__15636));
    LocalMux I__3477 (
            .O(N__15662),
            .I(N__15633));
    LocalMux I__3476 (
            .O(N__15659),
            .I(N__15630));
    LocalMux I__3475 (
            .O(N__15654),
            .I(N__15627));
    InMux I__3474 (
            .O(N__15653),
            .I(N__15620));
    InMux I__3473 (
            .O(N__15652),
            .I(N__15620));
    InMux I__3472 (
            .O(N__15651),
            .I(N__15620));
    LocalMux I__3471 (
            .O(N__15644),
            .I(N__15617));
    InMux I__3470 (
            .O(N__15643),
            .I(N__15612));
    InMux I__3469 (
            .O(N__15642),
            .I(N__15612));
    InMux I__3468 (
            .O(N__15641),
            .I(N__15605));
    InMux I__3467 (
            .O(N__15640),
            .I(N__15605));
    InMux I__3466 (
            .O(N__15639),
            .I(N__15605));
    Span4Mux_h I__3465 (
            .O(N__15636),
            .I(N__15598));
    Span4Mux_h I__3464 (
            .O(N__15633),
            .I(N__15598));
    Span4Mux_h I__3463 (
            .O(N__15630),
            .I(N__15598));
    Span4Mux_v I__3462 (
            .O(N__15627),
            .I(N__15591));
    LocalMux I__3461 (
            .O(N__15620),
            .I(N__15591));
    Span4Mux_s3_h I__3460 (
            .O(N__15617),
            .I(N__15591));
    LocalMux I__3459 (
            .O(N__15612),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3458 (
            .O(N__15605),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3457 (
            .O(N__15598),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3456 (
            .O(N__15591),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__3455 (
            .O(N__15582),
            .I(N__15574));
    InMux I__3454 (
            .O(N__15581),
            .I(N__15570));
    InMux I__3453 (
            .O(N__15580),
            .I(N__15567));
    CascadeMux I__3452 (
            .O(N__15579),
            .I(N__15564));
    InMux I__3451 (
            .O(N__15578),
            .I(N__15561));
    InMux I__3450 (
            .O(N__15577),
            .I(N__15557));
    LocalMux I__3449 (
            .O(N__15574),
            .I(N__15554));
    InMux I__3448 (
            .O(N__15573),
            .I(N__15551));
    LocalMux I__3447 (
            .O(N__15570),
            .I(N__15547));
    LocalMux I__3446 (
            .O(N__15567),
            .I(N__15544));
    InMux I__3445 (
            .O(N__15564),
            .I(N__15534));
    LocalMux I__3444 (
            .O(N__15561),
            .I(N__15531));
    InMux I__3443 (
            .O(N__15560),
            .I(N__15528));
    LocalMux I__3442 (
            .O(N__15557),
            .I(N__15521));
    Span4Mux_v I__3441 (
            .O(N__15554),
            .I(N__15521));
    LocalMux I__3440 (
            .O(N__15551),
            .I(N__15521));
    InMux I__3439 (
            .O(N__15550),
            .I(N__15518));
    Span4Mux_h I__3438 (
            .O(N__15547),
            .I(N__15515));
    Span4Mux_h I__3437 (
            .O(N__15544),
            .I(N__15512));
    InMux I__3436 (
            .O(N__15543),
            .I(N__15503));
    InMux I__3435 (
            .O(N__15542),
            .I(N__15503));
    InMux I__3434 (
            .O(N__15541),
            .I(N__15503));
    InMux I__3433 (
            .O(N__15540),
            .I(N__15503));
    InMux I__3432 (
            .O(N__15539),
            .I(N__15496));
    InMux I__3431 (
            .O(N__15538),
            .I(N__15496));
    InMux I__3430 (
            .O(N__15537),
            .I(N__15496));
    LocalMux I__3429 (
            .O(N__15534),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv12 I__3428 (
            .O(N__15531),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3427 (
            .O(N__15528),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__3426 (
            .O(N__15521),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3425 (
            .O(N__15518),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__3424 (
            .O(N__15515),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__3423 (
            .O(N__15512),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3422 (
            .O(N__15503),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3421 (
            .O(N__15496),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__3420 (
            .O(N__15477),
            .I(N__15467));
    InMux I__3419 (
            .O(N__15476),
            .I(N__15460));
    InMux I__3418 (
            .O(N__15475),
            .I(N__15460));
    InMux I__3417 (
            .O(N__15474),
            .I(N__15460));
    InMux I__3416 (
            .O(N__15473),
            .I(N__15453));
    InMux I__3415 (
            .O(N__15472),
            .I(N__15453));
    InMux I__3414 (
            .O(N__15471),
            .I(N__15453));
    InMux I__3413 (
            .O(N__15470),
            .I(N__15448));
    LocalMux I__3412 (
            .O(N__15467),
            .I(N__15445));
    LocalMux I__3411 (
            .O(N__15460),
            .I(N__15442));
    LocalMux I__3410 (
            .O(N__15453),
            .I(N__15439));
    InMux I__3409 (
            .O(N__15452),
            .I(N__15434));
    InMux I__3408 (
            .O(N__15451),
            .I(N__15434));
    LocalMux I__3407 (
            .O(N__15448),
            .I(N__15431));
    Span4Mux_v I__3406 (
            .O(N__15445),
            .I(N__15419));
    Span4Mux_s3_h I__3405 (
            .O(N__15442),
            .I(N__15419));
    Span4Mux_v I__3404 (
            .O(N__15439),
            .I(N__15419));
    LocalMux I__3403 (
            .O(N__15434),
            .I(N__15419));
    Span4Mux_h I__3402 (
            .O(N__15431),
            .I(N__15416));
    InMux I__3401 (
            .O(N__15430),
            .I(N__15411));
    InMux I__3400 (
            .O(N__15429),
            .I(N__15411));
    InMux I__3399 (
            .O(N__15428),
            .I(N__15408));
    Odrv4 I__3398 (
            .O(N__15419),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__3397 (
            .O(N__15416),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3396 (
            .O(N__15411),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3395 (
            .O(N__15408),
            .I(\uu2.un21_w_addr_displaying_i ));
    CascadeMux I__3394 (
            .O(N__15399),
            .I(N__15393));
    InMux I__3393 (
            .O(N__15398),
            .I(N__15390));
    CascadeMux I__3392 (
            .O(N__15397),
            .I(N__15387));
    InMux I__3391 (
            .O(N__15396),
            .I(N__15381));
    InMux I__3390 (
            .O(N__15393),
            .I(N__15381));
    LocalMux I__3389 (
            .O(N__15390),
            .I(N__15378));
    InMux I__3388 (
            .O(N__15387),
            .I(N__15375));
    CascadeMux I__3387 (
            .O(N__15386),
            .I(N__15370));
    LocalMux I__3386 (
            .O(N__15381),
            .I(N__15367));
    Span4Mux_v I__3385 (
            .O(N__15378),
            .I(N__15364));
    LocalMux I__3384 (
            .O(N__15375),
            .I(N__15361));
    InMux I__3383 (
            .O(N__15374),
            .I(N__15356));
    InMux I__3382 (
            .O(N__15373),
            .I(N__15356));
    InMux I__3381 (
            .O(N__15370),
            .I(N__15353));
    Span4Mux_v I__3380 (
            .O(N__15367),
            .I(N__15348));
    Span4Mux_h I__3379 (
            .O(N__15364),
            .I(N__15348));
    Odrv12 I__3378 (
            .O(N__15361),
            .I(\uu2.N_12_i ));
    LocalMux I__3377 (
            .O(N__15356),
            .I(\uu2.N_12_i ));
    LocalMux I__3376 (
            .O(N__15353),
            .I(\uu2.N_12_i ));
    Odrv4 I__3375 (
            .O(N__15348),
            .I(\uu2.N_12_i ));
    InMux I__3374 (
            .O(N__15339),
            .I(N__15336));
    LocalMux I__3373 (
            .O(N__15336),
            .I(N__15325));
    InMux I__3372 (
            .O(N__15335),
            .I(N__15322));
    InMux I__3371 (
            .O(N__15334),
            .I(N__15317));
    InMux I__3370 (
            .O(N__15333),
            .I(N__15317));
    InMux I__3369 (
            .O(N__15332),
            .I(N__15314));
    InMux I__3368 (
            .O(N__15331),
            .I(N__15306));
    InMux I__3367 (
            .O(N__15330),
            .I(N__15303));
    InMux I__3366 (
            .O(N__15329),
            .I(N__15300));
    InMux I__3365 (
            .O(N__15328),
            .I(N__15297));
    Span4Mux_h I__3364 (
            .O(N__15325),
            .I(N__15292));
    LocalMux I__3363 (
            .O(N__15322),
            .I(N__15292));
    LocalMux I__3362 (
            .O(N__15317),
            .I(N__15287));
    LocalMux I__3361 (
            .O(N__15314),
            .I(N__15287));
    InMux I__3360 (
            .O(N__15313),
            .I(N__15284));
    CascadeMux I__3359 (
            .O(N__15312),
            .I(N__15278));
    CascadeMux I__3358 (
            .O(N__15311),
            .I(N__15275));
    InMux I__3357 (
            .O(N__15310),
            .I(N__15270));
    InMux I__3356 (
            .O(N__15309),
            .I(N__15267));
    LocalMux I__3355 (
            .O(N__15306),
            .I(N__15262));
    LocalMux I__3354 (
            .O(N__15303),
            .I(N__15262));
    LocalMux I__3353 (
            .O(N__15300),
            .I(N__15256));
    LocalMux I__3352 (
            .O(N__15297),
            .I(N__15253));
    Span4Mux_h I__3351 (
            .O(N__15292),
            .I(N__15250));
    Span4Mux_h I__3350 (
            .O(N__15287),
            .I(N__15245));
    LocalMux I__3349 (
            .O(N__15284),
            .I(N__15245));
    InMux I__3348 (
            .O(N__15283),
            .I(N__15232));
    InMux I__3347 (
            .O(N__15282),
            .I(N__15232));
    InMux I__3346 (
            .O(N__15281),
            .I(N__15232));
    InMux I__3345 (
            .O(N__15278),
            .I(N__15232));
    InMux I__3344 (
            .O(N__15275),
            .I(N__15232));
    InMux I__3343 (
            .O(N__15274),
            .I(N__15232));
    InMux I__3342 (
            .O(N__15273),
            .I(N__15229));
    LocalMux I__3341 (
            .O(N__15270),
            .I(N__15222));
    LocalMux I__3340 (
            .O(N__15267),
            .I(N__15222));
    Span4Mux_h I__3339 (
            .O(N__15262),
            .I(N__15222));
    InMux I__3338 (
            .O(N__15261),
            .I(N__15215));
    InMux I__3337 (
            .O(N__15260),
            .I(N__15215));
    InMux I__3336 (
            .O(N__15259),
            .I(N__15215));
    Odrv4 I__3335 (
            .O(N__15256),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__3334 (
            .O(N__15253),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__3333 (
            .O(N__15250),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__3332 (
            .O(N__15245),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__3331 (
            .O(N__15232),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__3330 (
            .O(N__15229),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__3329 (
            .O(N__15222),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__3328 (
            .O(N__15215),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__3327 (
            .O(N__15198),
            .I(N__15193));
    InMux I__3326 (
            .O(N__15197),
            .I(N__15184));
    CascadeMux I__3325 (
            .O(N__15196),
            .I(N__15180));
    LocalMux I__3324 (
            .O(N__15193),
            .I(N__15176));
    InMux I__3323 (
            .O(N__15192),
            .I(N__15173));
    InMux I__3322 (
            .O(N__15191),
            .I(N__15170));
    CascadeMux I__3321 (
            .O(N__15190),
            .I(N__15167));
    InMux I__3320 (
            .O(N__15189),
            .I(N__15162));
    InMux I__3319 (
            .O(N__15188),
            .I(N__15162));
    InMux I__3318 (
            .O(N__15187),
            .I(N__15159));
    LocalMux I__3317 (
            .O(N__15184),
            .I(N__15153));
    InMux I__3316 (
            .O(N__15183),
            .I(N__15150));
    InMux I__3315 (
            .O(N__15180),
            .I(N__15144));
    InMux I__3314 (
            .O(N__15179),
            .I(N__15144));
    Span4Mux_h I__3313 (
            .O(N__15176),
            .I(N__15139));
    LocalMux I__3312 (
            .O(N__15173),
            .I(N__15139));
    LocalMux I__3311 (
            .O(N__15170),
            .I(N__15136));
    InMux I__3310 (
            .O(N__15167),
            .I(N__15133));
    LocalMux I__3309 (
            .O(N__15162),
            .I(N__15128));
    LocalMux I__3308 (
            .O(N__15159),
            .I(N__15128));
    CascadeMux I__3307 (
            .O(N__15158),
            .I(N__15125));
    InMux I__3306 (
            .O(N__15157),
            .I(N__15119));
    InMux I__3305 (
            .O(N__15156),
            .I(N__15119));
    Span4Mux_h I__3304 (
            .O(N__15153),
            .I(N__15114));
    LocalMux I__3303 (
            .O(N__15150),
            .I(N__15114));
    InMux I__3302 (
            .O(N__15149),
            .I(N__15107));
    LocalMux I__3301 (
            .O(N__15144),
            .I(N__15104));
    Span4Mux_h I__3300 (
            .O(N__15139),
            .I(N__15101));
    Span4Mux_h I__3299 (
            .O(N__15136),
            .I(N__15098));
    LocalMux I__3298 (
            .O(N__15133),
            .I(N__15093));
    Span4Mux_h I__3297 (
            .O(N__15128),
            .I(N__15093));
    InMux I__3296 (
            .O(N__15125),
            .I(N__15090));
    InMux I__3295 (
            .O(N__15124),
            .I(N__15087));
    LocalMux I__3294 (
            .O(N__15119),
            .I(N__15082));
    Span4Mux_h I__3293 (
            .O(N__15114),
            .I(N__15082));
    InMux I__3292 (
            .O(N__15113),
            .I(N__15073));
    InMux I__3291 (
            .O(N__15112),
            .I(N__15073));
    InMux I__3290 (
            .O(N__15111),
            .I(N__15073));
    InMux I__3289 (
            .O(N__15110),
            .I(N__15073));
    LocalMux I__3288 (
            .O(N__15107),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3287 (
            .O(N__15104),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3286 (
            .O(N__15101),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3285 (
            .O(N__15098),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3284 (
            .O(N__15093),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3283 (
            .O(N__15090),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3282 (
            .O(N__15087),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3281 (
            .O(N__15082),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3280 (
            .O(N__15073),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__3279 (
            .O(N__15054),
            .I(N__15045));
    InMux I__3278 (
            .O(N__15053),
            .I(N__15045));
    InMux I__3277 (
            .O(N__15052),
            .I(N__15040));
    InMux I__3276 (
            .O(N__15051),
            .I(N__15035));
    InMux I__3275 (
            .O(N__15050),
            .I(N__15035));
    LocalMux I__3274 (
            .O(N__15045),
            .I(N__15032));
    InMux I__3273 (
            .O(N__15044),
            .I(N__15029));
    InMux I__3272 (
            .O(N__15043),
            .I(N__15026));
    LocalMux I__3271 (
            .O(N__15040),
            .I(N__15023));
    LocalMux I__3270 (
            .O(N__15035),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__3269 (
            .O(N__15032),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3268 (
            .O(N__15029),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3267 (
            .O(N__15026),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv12 I__3266 (
            .O(N__15023),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    CascadeMux I__3265 (
            .O(N__15012),
            .I(\uu2.N_272_cascade_ ));
    InMux I__3264 (
            .O(N__15009),
            .I(N__15006));
    LocalMux I__3263 (
            .O(N__15006),
            .I(\uu2.mem0.m317_0_a6_1_0 ));
    InMux I__3262 (
            .O(N__15003),
            .I(N__15000));
    LocalMux I__3261 (
            .O(N__15000),
            .I(\uu2.mem0.N_13 ));
    InMux I__3260 (
            .O(N__14997),
            .I(N__14994));
    LocalMux I__3259 (
            .O(N__14994),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__3258 (
            .O(N__14991),
            .I(N__14967));
    InMux I__3257 (
            .O(N__14990),
            .I(N__14967));
    InMux I__3256 (
            .O(N__14989),
            .I(N__14967));
    InMux I__3255 (
            .O(N__14988),
            .I(N__14960));
    InMux I__3254 (
            .O(N__14987),
            .I(N__14960));
    InMux I__3253 (
            .O(N__14986),
            .I(N__14960));
    InMux I__3252 (
            .O(N__14985),
            .I(N__14953));
    InMux I__3251 (
            .O(N__14984),
            .I(N__14953));
    InMux I__3250 (
            .O(N__14983),
            .I(N__14953));
    InMux I__3249 (
            .O(N__14982),
            .I(N__14942));
    InMux I__3248 (
            .O(N__14981),
            .I(N__14942));
    InMux I__3247 (
            .O(N__14980),
            .I(N__14937));
    InMux I__3246 (
            .O(N__14979),
            .I(N__14937));
    InMux I__3245 (
            .O(N__14978),
            .I(N__14927));
    InMux I__3244 (
            .O(N__14977),
            .I(N__14927));
    InMux I__3243 (
            .O(N__14976),
            .I(N__14927));
    InMux I__3242 (
            .O(N__14975),
            .I(N__14922));
    InMux I__3241 (
            .O(N__14974),
            .I(N__14922));
    LocalMux I__3240 (
            .O(N__14967),
            .I(N__14919));
    LocalMux I__3239 (
            .O(N__14960),
            .I(N__14914));
    LocalMux I__3238 (
            .O(N__14953),
            .I(N__14914));
    InMux I__3237 (
            .O(N__14952),
            .I(N__14903));
    InMux I__3236 (
            .O(N__14951),
            .I(N__14903));
    InMux I__3235 (
            .O(N__14950),
            .I(N__14903));
    InMux I__3234 (
            .O(N__14949),
            .I(N__14903));
    InMux I__3233 (
            .O(N__14948),
            .I(N__14903));
    InMux I__3232 (
            .O(N__14947),
            .I(N__14897));
    LocalMux I__3231 (
            .O(N__14942),
            .I(N__14892));
    LocalMux I__3230 (
            .O(N__14937),
            .I(N__14892));
    InMux I__3229 (
            .O(N__14936),
            .I(N__14887));
    InMux I__3228 (
            .O(N__14935),
            .I(N__14887));
    CascadeMux I__3227 (
            .O(N__14934),
            .I(N__14883));
    LocalMux I__3226 (
            .O(N__14927),
            .I(N__14878));
    LocalMux I__3225 (
            .O(N__14922),
            .I(N__14878));
    Span4Mux_s3_v I__3224 (
            .O(N__14919),
            .I(N__14873));
    Span4Mux_h I__3223 (
            .O(N__14914),
            .I(N__14873));
    LocalMux I__3222 (
            .O(N__14903),
            .I(N__14870));
    InMux I__3221 (
            .O(N__14902),
            .I(N__14863));
    InMux I__3220 (
            .O(N__14901),
            .I(N__14863));
    InMux I__3219 (
            .O(N__14900),
            .I(N__14863));
    LocalMux I__3218 (
            .O(N__14897),
            .I(N__14860));
    Span4Mux_v I__3217 (
            .O(N__14892),
            .I(N__14855));
    LocalMux I__3216 (
            .O(N__14887),
            .I(N__14855));
    InMux I__3215 (
            .O(N__14886),
            .I(N__14850));
    InMux I__3214 (
            .O(N__14883),
            .I(N__14850));
    Span12Mux_s10_v I__3213 (
            .O(N__14878),
            .I(N__14847));
    Span4Mux_v I__3212 (
            .O(N__14873),
            .I(N__14840));
    Span4Mux_h I__3211 (
            .O(N__14870),
            .I(N__14840));
    LocalMux I__3210 (
            .O(N__14863),
            .I(N__14840));
    Span4Mux_h I__3209 (
            .O(N__14860),
            .I(N__14837));
    Span4Mux_v I__3208 (
            .O(N__14855),
            .I(N__14832));
    LocalMux I__3207 (
            .O(N__14850),
            .I(N__14832));
    Odrv12 I__3206 (
            .O(N__14847),
            .I(\Lab_UT.Run ));
    Odrv4 I__3205 (
            .O(N__14840),
            .I(\Lab_UT.Run ));
    Odrv4 I__3204 (
            .O(N__14837),
            .I(\Lab_UT.Run ));
    Odrv4 I__3203 (
            .O(N__14832),
            .I(\Lab_UT.Run ));
    InMux I__3202 (
            .O(N__14823),
            .I(N__14820));
    LocalMux I__3201 (
            .O(N__14820),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__3200 (
            .O(N__14817),
            .I(N__14811));
    InMux I__3199 (
            .O(N__14816),
            .I(N__14811));
    LocalMux I__3198 (
            .O(N__14811),
            .I(N__14808));
    Odrv12 I__3197 (
            .O(N__14808),
            .I(\uu2.bitmapZ0Z_314 ));
    CascadeMux I__3196 (
            .O(N__14805),
            .I(N__14799));
    InMux I__3195 (
            .O(N__14804),
            .I(N__14794));
    InMux I__3194 (
            .O(N__14803),
            .I(N__14794));
    InMux I__3193 (
            .O(N__14802),
            .I(N__14790));
    InMux I__3192 (
            .O(N__14799),
            .I(N__14787));
    LocalMux I__3191 (
            .O(N__14794),
            .I(N__14781));
    InMux I__3190 (
            .O(N__14793),
            .I(N__14778));
    LocalMux I__3189 (
            .O(N__14790),
            .I(N__14775));
    LocalMux I__3188 (
            .O(N__14787),
            .I(N__14772));
    InMux I__3187 (
            .O(N__14786),
            .I(N__14769));
    InMux I__3186 (
            .O(N__14785),
            .I(N__14766));
    InMux I__3185 (
            .O(N__14784),
            .I(N__14763));
    Span4Mux_h I__3184 (
            .O(N__14781),
            .I(N__14758));
    LocalMux I__3183 (
            .O(N__14778),
            .I(N__14758));
    Span4Mux_v I__3182 (
            .O(N__14775),
            .I(N__14753));
    Span4Mux_v I__3181 (
            .O(N__14772),
            .I(N__14753));
    LocalMux I__3180 (
            .O(N__14769),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__3179 (
            .O(N__14766),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__3178 (
            .O(N__14763),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    Odrv4 I__3177 (
            .O(N__14758),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    Odrv4 I__3176 (
            .O(N__14753),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    InMux I__3175 (
            .O(N__14742),
            .I(N__14739));
    LocalMux I__3174 (
            .O(N__14739),
            .I(\uu2.N_272 ));
    InMux I__3173 (
            .O(N__14736),
            .I(N__14733));
    LocalMux I__3172 (
            .O(N__14733),
            .I(N__14728));
    InMux I__3171 (
            .O(N__14732),
            .I(N__14725));
    InMux I__3170 (
            .O(N__14731),
            .I(N__14722));
    Span4Mux_v I__3169 (
            .O(N__14728),
            .I(N__14717));
    LocalMux I__3168 (
            .O(N__14725),
            .I(N__14717));
    LocalMux I__3167 (
            .O(N__14722),
            .I(N__14714));
    Span4Mux_h I__3166 (
            .O(N__14717),
            .I(N__14711));
    Span12Mux_s10_h I__3165 (
            .O(N__14714),
            .I(N__14708));
    Span4Mux_s2_h I__3164 (
            .O(N__14711),
            .I(N__14705));
    Odrv12 I__3163 (
            .O(N__14708),
            .I(\uu2.bitmapZ0Z_111 ));
    Odrv4 I__3162 (
            .O(N__14705),
            .I(\uu2.bitmapZ0Z_111 ));
    CascadeMux I__3161 (
            .O(N__14700),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_ ));
    InMux I__3160 (
            .O(N__14697),
            .I(N__14694));
    LocalMux I__3159 (
            .O(N__14694),
            .I(\uu2.mem0.bitmap_pmux_u_i_4_0 ));
    InMux I__3158 (
            .O(N__14691),
            .I(N__14688));
    LocalMux I__3157 (
            .O(N__14688),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_69 ));
    InMux I__3156 (
            .O(N__14685),
            .I(N__14677));
    InMux I__3155 (
            .O(N__14684),
            .I(N__14677));
    CascadeMux I__3154 (
            .O(N__14683),
            .I(N__14674));
    InMux I__3153 (
            .O(N__14682),
            .I(N__14671));
    LocalMux I__3152 (
            .O(N__14677),
            .I(N__14665));
    InMux I__3151 (
            .O(N__14674),
            .I(N__14662));
    LocalMux I__3150 (
            .O(N__14671),
            .I(N__14659));
    CascadeMux I__3149 (
            .O(N__14670),
            .I(N__14656));
    CascadeMux I__3148 (
            .O(N__14669),
            .I(N__14653));
    InMux I__3147 (
            .O(N__14668),
            .I(N__14646));
    Span4Mux_v I__3146 (
            .O(N__14665),
            .I(N__14641));
    LocalMux I__3145 (
            .O(N__14662),
            .I(N__14641));
    Span4Mux_v I__3144 (
            .O(N__14659),
            .I(N__14638));
    InMux I__3143 (
            .O(N__14656),
            .I(N__14635));
    InMux I__3142 (
            .O(N__14653),
            .I(N__14632));
    InMux I__3141 (
            .O(N__14652),
            .I(N__14629));
    CascadeMux I__3140 (
            .O(N__14651),
            .I(N__14626));
    CascadeMux I__3139 (
            .O(N__14650),
            .I(N__14622));
    CascadeMux I__3138 (
            .O(N__14649),
            .I(N__14617));
    LocalMux I__3137 (
            .O(N__14646),
            .I(N__14614));
    Span4Mux_h I__3136 (
            .O(N__14641),
            .I(N__14611));
    Span4Mux_h I__3135 (
            .O(N__14638),
            .I(N__14602));
    LocalMux I__3134 (
            .O(N__14635),
            .I(N__14602));
    LocalMux I__3133 (
            .O(N__14632),
            .I(N__14602));
    LocalMux I__3132 (
            .O(N__14629),
            .I(N__14602));
    InMux I__3131 (
            .O(N__14626),
            .I(N__14589));
    InMux I__3130 (
            .O(N__14625),
            .I(N__14589));
    InMux I__3129 (
            .O(N__14622),
            .I(N__14589));
    InMux I__3128 (
            .O(N__14621),
            .I(N__14589));
    InMux I__3127 (
            .O(N__14620),
            .I(N__14589));
    InMux I__3126 (
            .O(N__14617),
            .I(N__14589));
    Odrv12 I__3125 (
            .O(N__14614),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__3124 (
            .O(N__14611),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__3123 (
            .O(N__14602),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3122 (
            .O(N__14589),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CEMux I__3121 (
            .O(N__14580),
            .I(N__14575));
    CEMux I__3120 (
            .O(N__14579),
            .I(N__14572));
    CEMux I__3119 (
            .O(N__14578),
            .I(N__14569));
    LocalMux I__3118 (
            .O(N__14575),
            .I(N__14566));
    LocalMux I__3117 (
            .O(N__14572),
            .I(N__14563));
    LocalMux I__3116 (
            .O(N__14569),
            .I(N__14560));
    Span4Mux_h I__3115 (
            .O(N__14566),
            .I(N__14557));
    Span4Mux_v I__3114 (
            .O(N__14563),
            .I(N__14554));
    Span4Mux_v I__3113 (
            .O(N__14560),
            .I(N__14551));
    Odrv4 I__3112 (
            .O(N__14557),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    Odrv4 I__3111 (
            .O(N__14554),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    Odrv4 I__3110 (
            .O(N__14551),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    CascadeMux I__3109 (
            .O(N__14544),
            .I(\uu2.mem0.G_13_0_a2_1_cascade_ ));
    InMux I__3108 (
            .O(N__14541),
            .I(N__14538));
    LocalMux I__3107 (
            .O(N__14538),
            .I(N__14535));
    Odrv12 I__3106 (
            .O(N__14535),
            .I(\uu2.mem0.G_13_0_a3_1_2 ));
    CascadeMux I__3105 (
            .O(N__14532),
            .I(N__14522));
    InMux I__3104 (
            .O(N__14531),
            .I(N__14516));
    InMux I__3103 (
            .O(N__14530),
            .I(N__14513));
    InMux I__3102 (
            .O(N__14529),
            .I(N__14510));
    InMux I__3101 (
            .O(N__14528),
            .I(N__14505));
    InMux I__3100 (
            .O(N__14527),
            .I(N__14505));
    InMux I__3099 (
            .O(N__14526),
            .I(N__14498));
    InMux I__3098 (
            .O(N__14525),
            .I(N__14498));
    InMux I__3097 (
            .O(N__14522),
            .I(N__14493));
    InMux I__3096 (
            .O(N__14521),
            .I(N__14493));
    InMux I__3095 (
            .O(N__14520),
            .I(N__14488));
    InMux I__3094 (
            .O(N__14519),
            .I(N__14488));
    LocalMux I__3093 (
            .O(N__14516),
            .I(N__14481));
    LocalMux I__3092 (
            .O(N__14513),
            .I(N__14481));
    LocalMux I__3091 (
            .O(N__14510),
            .I(N__14478));
    LocalMux I__3090 (
            .O(N__14505),
            .I(N__14475));
    InMux I__3089 (
            .O(N__14504),
            .I(N__14470));
    InMux I__3088 (
            .O(N__14503),
            .I(N__14470));
    LocalMux I__3087 (
            .O(N__14498),
            .I(N__14463));
    LocalMux I__3086 (
            .O(N__14493),
            .I(N__14463));
    LocalMux I__3085 (
            .O(N__14488),
            .I(N__14463));
    InMux I__3084 (
            .O(N__14487),
            .I(N__14457));
    InMux I__3083 (
            .O(N__14486),
            .I(N__14454));
    Span4Mux_v I__3082 (
            .O(N__14481),
            .I(N__14451));
    Span4Mux_v I__3081 (
            .O(N__14478),
            .I(N__14442));
    Span4Mux_v I__3080 (
            .O(N__14475),
            .I(N__14442));
    LocalMux I__3079 (
            .O(N__14470),
            .I(N__14442));
    Span4Mux_h I__3078 (
            .O(N__14463),
            .I(N__14442));
    InMux I__3077 (
            .O(N__14462),
            .I(N__14437));
    InMux I__3076 (
            .O(N__14461),
            .I(N__14437));
    InMux I__3075 (
            .O(N__14460),
            .I(N__14434));
    LocalMux I__3074 (
            .O(N__14457),
            .I(L3_tx_data_rdy));
    LocalMux I__3073 (
            .O(N__14454),
            .I(L3_tx_data_rdy));
    Odrv4 I__3072 (
            .O(N__14451),
            .I(L3_tx_data_rdy));
    Odrv4 I__3071 (
            .O(N__14442),
            .I(L3_tx_data_rdy));
    LocalMux I__3070 (
            .O(N__14437),
            .I(L3_tx_data_rdy));
    LocalMux I__3069 (
            .O(N__14434),
            .I(L3_tx_data_rdy));
    InMux I__3068 (
            .O(N__14421),
            .I(N__14418));
    LocalMux I__3067 (
            .O(N__14418),
            .I(N__14415));
    Span4Mux_h I__3066 (
            .O(N__14415),
            .I(N__14410));
    InMux I__3065 (
            .O(N__14414),
            .I(N__14405));
    InMux I__3064 (
            .O(N__14413),
            .I(N__14405));
    Odrv4 I__3063 (
            .O(N__14410),
            .I(L3_tx_data_1));
    LocalMux I__3062 (
            .O(N__14405),
            .I(L3_tx_data_1));
    CascadeMux I__3061 (
            .O(N__14400),
            .I(\uu2.mem0.G_13_0_a2_2_cascade_ ));
    CascadeMux I__3060 (
            .O(N__14397),
            .I(N__14391));
    InMux I__3059 (
            .O(N__14396),
            .I(N__14381));
    InMux I__3058 (
            .O(N__14395),
            .I(N__14376));
    InMux I__3057 (
            .O(N__14394),
            .I(N__14376));
    InMux I__3056 (
            .O(N__14391),
            .I(N__14371));
    InMux I__3055 (
            .O(N__14390),
            .I(N__14362));
    InMux I__3054 (
            .O(N__14389),
            .I(N__14362));
    InMux I__3053 (
            .O(N__14388),
            .I(N__14362));
    InMux I__3052 (
            .O(N__14387),
            .I(N__14362));
    InMux I__3051 (
            .O(N__14386),
            .I(N__14357));
    InMux I__3050 (
            .O(N__14385),
            .I(N__14357));
    InMux I__3049 (
            .O(N__14384),
            .I(N__14354));
    LocalMux I__3048 (
            .O(N__14381),
            .I(N__14348));
    LocalMux I__3047 (
            .O(N__14376),
            .I(N__14345));
    InMux I__3046 (
            .O(N__14375),
            .I(N__14340));
    InMux I__3045 (
            .O(N__14374),
            .I(N__14340));
    LocalMux I__3044 (
            .O(N__14371),
            .I(N__14337));
    LocalMux I__3043 (
            .O(N__14362),
            .I(N__14332));
    LocalMux I__3042 (
            .O(N__14357),
            .I(N__14332));
    LocalMux I__3041 (
            .O(N__14354),
            .I(N__14329));
    InMux I__3040 (
            .O(N__14353),
            .I(N__14325));
    InMux I__3039 (
            .O(N__14352),
            .I(N__14320));
    InMux I__3038 (
            .O(N__14351),
            .I(N__14320));
    Span4Mux_v I__3037 (
            .O(N__14348),
            .I(N__14313));
    Span4Mux_h I__3036 (
            .O(N__14345),
            .I(N__14313));
    LocalMux I__3035 (
            .O(N__14340),
            .I(N__14313));
    Span4Mux_h I__3034 (
            .O(N__14337),
            .I(N__14308));
    Span4Mux_h I__3033 (
            .O(N__14332),
            .I(N__14308));
    Span4Mux_h I__3032 (
            .O(N__14329),
            .I(N__14305));
    InMux I__3031 (
            .O(N__14328),
            .I(N__14302));
    LocalMux I__3030 (
            .O(N__14325),
            .I(N_96));
    LocalMux I__3029 (
            .O(N__14320),
            .I(N_96));
    Odrv4 I__3028 (
            .O(N__14313),
            .I(N_96));
    Odrv4 I__3027 (
            .O(N__14308),
            .I(N_96));
    Odrv4 I__3026 (
            .O(N__14305),
            .I(N_96));
    LocalMux I__3025 (
            .O(N__14302),
            .I(N_96));
    InMux I__3024 (
            .O(N__14289),
            .I(N__14286));
    LocalMux I__3023 (
            .O(N__14286),
            .I(N__14283));
    Span4Mux_h I__3022 (
            .O(N__14283),
            .I(N__14280));
    Odrv4 I__3021 (
            .O(N__14280),
            .I(\uu2.mem0.G_13_0_0 ));
    InMux I__3020 (
            .O(N__14277),
            .I(N__14274));
    LocalMux I__3019 (
            .O(N__14274),
            .I(N__14271));
    Odrv4 I__3018 (
            .O(N__14271),
            .I(\uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0 ));
    InMux I__3017 (
            .O(N__14268),
            .I(N__14261));
    InMux I__3016 (
            .O(N__14267),
            .I(N__14261));
    InMux I__3015 (
            .O(N__14266),
            .I(N__14256));
    LocalMux I__3014 (
            .O(N__14261),
            .I(N__14252));
    InMux I__3013 (
            .O(N__14260),
            .I(N__14247));
    InMux I__3012 (
            .O(N__14259),
            .I(N__14247));
    LocalMux I__3011 (
            .O(N__14256),
            .I(N__14238));
    InMux I__3010 (
            .O(N__14255),
            .I(N__14235));
    Span4Mux_h I__3009 (
            .O(N__14252),
            .I(N__14232));
    LocalMux I__3008 (
            .O(N__14247),
            .I(N__14229));
    InMux I__3007 (
            .O(N__14246),
            .I(N__14224));
    InMux I__3006 (
            .O(N__14245),
            .I(N__14224));
    InMux I__3005 (
            .O(N__14244),
            .I(N__14217));
    InMux I__3004 (
            .O(N__14243),
            .I(N__14217));
    InMux I__3003 (
            .O(N__14242),
            .I(N__14217));
    InMux I__3002 (
            .O(N__14241),
            .I(N__14213));
    Span4Mux_v I__3001 (
            .O(N__14238),
            .I(N__14208));
    LocalMux I__3000 (
            .O(N__14235),
            .I(N__14208));
    Span4Mux_v I__2999 (
            .O(N__14232),
            .I(N__14205));
    Span4Mux_v I__2998 (
            .O(N__14229),
            .I(N__14202));
    LocalMux I__2997 (
            .O(N__14224),
            .I(N__14197));
    LocalMux I__2996 (
            .O(N__14217),
            .I(N__14197));
    InMux I__2995 (
            .O(N__14216),
            .I(N__14194));
    LocalMux I__2994 (
            .O(N__14213),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__2993 (
            .O(N__14208),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__2992 (
            .O(N__14205),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__2991 (
            .O(N__14202),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv12 I__2990 (
            .O(N__14197),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__2989 (
            .O(N__14194),
            .I(\Lab_UT.di_Mones_0 ));
    InMux I__2988 (
            .O(N__14181),
            .I(N__14172));
    InMux I__2987 (
            .O(N__14180),
            .I(N__14172));
    InMux I__2986 (
            .O(N__14179),
            .I(N__14167));
    InMux I__2985 (
            .O(N__14178),
            .I(N__14167));
    InMux I__2984 (
            .O(N__14177),
            .I(N__14163));
    LocalMux I__2983 (
            .O(N__14172),
            .I(N__14155));
    LocalMux I__2982 (
            .O(N__14167),
            .I(N__14155));
    InMux I__2981 (
            .O(N__14166),
            .I(N__14151));
    LocalMux I__2980 (
            .O(N__14163),
            .I(N__14148));
    InMux I__2979 (
            .O(N__14162),
            .I(N__14143));
    InMux I__2978 (
            .O(N__14161),
            .I(N__14143));
    InMux I__2977 (
            .O(N__14160),
            .I(N__14140));
    Span4Mux_h I__2976 (
            .O(N__14155),
            .I(N__14137));
    InMux I__2975 (
            .O(N__14154),
            .I(N__14133));
    LocalMux I__2974 (
            .O(N__14151),
            .I(N__14130));
    Span4Mux_h I__2973 (
            .O(N__14148),
            .I(N__14125));
    LocalMux I__2972 (
            .O(N__14143),
            .I(N__14125));
    LocalMux I__2971 (
            .O(N__14140),
            .I(N__14120));
    Span4Mux_v I__2970 (
            .O(N__14137),
            .I(N__14120));
    InMux I__2969 (
            .O(N__14136),
            .I(N__14117));
    LocalMux I__2968 (
            .O(N__14133),
            .I(N__14114));
    Odrv4 I__2967 (
            .O(N__14130),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__2966 (
            .O(N__14125),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__2965 (
            .O(N__14120),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__2964 (
            .O(N__14117),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv12 I__2963 (
            .O(N__14114),
            .I(\Lab_UT.di_Mones_3 ));
    InMux I__2962 (
            .O(N__14103),
            .I(N__14095));
    InMux I__2961 (
            .O(N__14102),
            .I(N__14092));
    CascadeMux I__2960 (
            .O(N__14101),
            .I(N__14089));
    CascadeMux I__2959 (
            .O(N__14100),
            .I(N__14086));
    CascadeMux I__2958 (
            .O(N__14099),
            .I(N__14080));
    CascadeMux I__2957 (
            .O(N__14098),
            .I(N__14077));
    LocalMux I__2956 (
            .O(N__14095),
            .I(N__14073));
    LocalMux I__2955 (
            .O(N__14092),
            .I(N__14070));
    InMux I__2954 (
            .O(N__14089),
            .I(N__14065));
    InMux I__2953 (
            .O(N__14086),
            .I(N__14065));
    CascadeMux I__2952 (
            .O(N__14085),
            .I(N__14062));
    CascadeMux I__2951 (
            .O(N__14084),
            .I(N__14059));
    CascadeMux I__2950 (
            .O(N__14083),
            .I(N__14054));
    InMux I__2949 (
            .O(N__14080),
            .I(N__14049));
    InMux I__2948 (
            .O(N__14077),
            .I(N__14049));
    InMux I__2947 (
            .O(N__14076),
            .I(N__14046));
    Span4Mux_v I__2946 (
            .O(N__14073),
            .I(N__14043));
    Span12Mux_v I__2945 (
            .O(N__14070),
            .I(N__14038));
    LocalMux I__2944 (
            .O(N__14065),
            .I(N__14038));
    InMux I__2943 (
            .O(N__14062),
            .I(N__14033));
    InMux I__2942 (
            .O(N__14059),
            .I(N__14033));
    InMux I__2941 (
            .O(N__14058),
            .I(N__14026));
    InMux I__2940 (
            .O(N__14057),
            .I(N__14026));
    InMux I__2939 (
            .O(N__14054),
            .I(N__14026));
    LocalMux I__2938 (
            .O(N__14049),
            .I(N__14021));
    LocalMux I__2937 (
            .O(N__14046),
            .I(N__14021));
    Odrv4 I__2936 (
            .O(N__14043),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv12 I__2935 (
            .O(N__14038),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2934 (
            .O(N__14033),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2933 (
            .O(N__14026),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv12 I__2932 (
            .O(N__14021),
            .I(\Lab_UT.di_Mones_1 ));
    CascadeMux I__2931 (
            .O(N__14010),
            .I(\Lab_UT.bcd2segment1.N_248_cascade_ ));
    InMux I__2930 (
            .O(N__14007),
            .I(N__14004));
    LocalMux I__2929 (
            .O(N__14004),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__2928 (
            .O(N__14001),
            .I(N__13998));
    LocalMux I__2927 (
            .O(N__13998),
            .I(\uu2.bitmapZ0Z_72 ));
    InMux I__2926 (
            .O(N__13995),
            .I(N__13992));
    LocalMux I__2925 (
            .O(N__13992),
            .I(\uu2.m76_bm_1_0 ));
    InMux I__2924 (
            .O(N__13989),
            .I(N__13986));
    LocalMux I__2923 (
            .O(N__13986),
            .I(N__13982));
    CascadeMux I__2922 (
            .O(N__13985),
            .I(N__13977));
    Span4Mux_h I__2921 (
            .O(N__13982),
            .I(N__13974));
    InMux I__2920 (
            .O(N__13981),
            .I(N__13971));
    InMux I__2919 (
            .O(N__13980),
            .I(N__13966));
    InMux I__2918 (
            .O(N__13977),
            .I(N__13966));
    Odrv4 I__2917 (
            .O(N__13974),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__2916 (
            .O(N__13971),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__2915 (
            .O(N__13966),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__2914 (
            .O(N__13959),
            .I(N__13956));
    LocalMux I__2913 (
            .O(N__13956),
            .I(N__13953));
    Span4Mux_h I__2912 (
            .O(N__13953),
            .I(N__13950));
    Span4Mux_h I__2911 (
            .O(N__13950),
            .I(N__13947));
    Odrv4 I__2910 (
            .O(N__13947),
            .I(\uu2.mem0.g1_2_2 ));
    InMux I__2909 (
            .O(N__13944),
            .I(N__13941));
    LocalMux I__2908 (
            .O(N__13941),
            .I(N__13938));
    Span12Mux_s8_h I__2907 (
            .O(N__13938),
            .I(N__13935));
    Odrv12 I__2906 (
            .O(N__13935),
            .I(\uu2.mem0.g2_0_0_0_0 ));
    InMux I__2905 (
            .O(N__13932),
            .I(N__13929));
    LocalMux I__2904 (
            .O(N__13929),
            .I(N__13926));
    Span4Mux_h I__2903 (
            .O(N__13926),
            .I(N__13923));
    Odrv4 I__2902 (
            .O(N__13923),
            .I(\uu2.mem0.g2_2 ));
    CascadeMux I__2901 (
            .O(N__13920),
            .I(N__13914));
    CascadeMux I__2900 (
            .O(N__13919),
            .I(N__13909));
    CascadeMux I__2899 (
            .O(N__13918),
            .I(N__13905));
    CascadeMux I__2898 (
            .O(N__13917),
            .I(N__13901));
    InMux I__2897 (
            .O(N__13914),
            .I(N__13897));
    InMux I__2896 (
            .O(N__13913),
            .I(N__13894));
    InMux I__2895 (
            .O(N__13912),
            .I(N__13891));
    InMux I__2894 (
            .O(N__13909),
            .I(N__13888));
    InMux I__2893 (
            .O(N__13908),
            .I(N__13884));
    InMux I__2892 (
            .O(N__13905),
            .I(N__13881));
    InMux I__2891 (
            .O(N__13904),
            .I(N__13874));
    InMux I__2890 (
            .O(N__13901),
            .I(N__13874));
    InMux I__2889 (
            .O(N__13900),
            .I(N__13874));
    LocalMux I__2888 (
            .O(N__13897),
            .I(N__13871));
    LocalMux I__2887 (
            .O(N__13894),
            .I(N__13868));
    LocalMux I__2886 (
            .O(N__13891),
            .I(N__13865));
    LocalMux I__2885 (
            .O(N__13888),
            .I(N__13862));
    InMux I__2884 (
            .O(N__13887),
            .I(N__13859));
    LocalMux I__2883 (
            .O(N__13884),
            .I(N__13856));
    LocalMux I__2882 (
            .O(N__13881),
            .I(N__13851));
    LocalMux I__2881 (
            .O(N__13874),
            .I(N__13851));
    Span4Mux_v I__2880 (
            .O(N__13871),
            .I(N__13842));
    Span4Mux_h I__2879 (
            .O(N__13868),
            .I(N__13842));
    Span4Mux_h I__2878 (
            .O(N__13865),
            .I(N__13842));
    Span4Mux_h I__2877 (
            .O(N__13862),
            .I(N__13842));
    LocalMux I__2876 (
            .O(N__13859),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__2875 (
            .O(N__13856),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__2874 (
            .O(N__13851),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__2873 (
            .O(N__13842),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    InMux I__2872 (
            .O(N__13833),
            .I(N__13830));
    LocalMux I__2871 (
            .O(N__13830),
            .I(N__13823));
    InMux I__2870 (
            .O(N__13829),
            .I(N__13820));
    CascadeMux I__2869 (
            .O(N__13828),
            .I(N__13817));
    CascadeMux I__2868 (
            .O(N__13827),
            .I(N__13812));
    InMux I__2867 (
            .O(N__13826),
            .I(N__13807));
    Span4Mux_h I__2866 (
            .O(N__13823),
            .I(N__13804));
    LocalMux I__2865 (
            .O(N__13820),
            .I(N__13801));
    InMux I__2864 (
            .O(N__13817),
            .I(N__13794));
    InMux I__2863 (
            .O(N__13816),
            .I(N__13794));
    InMux I__2862 (
            .O(N__13815),
            .I(N__13794));
    InMux I__2861 (
            .O(N__13812),
            .I(N__13787));
    InMux I__2860 (
            .O(N__13811),
            .I(N__13787));
    InMux I__2859 (
            .O(N__13810),
            .I(N__13787));
    LocalMux I__2858 (
            .O(N__13807),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv4 I__2857 (
            .O(N__13804),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv12 I__2856 (
            .O(N__13801),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2855 (
            .O(N__13794),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2854 (
            .O(N__13787),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    InMux I__2853 (
            .O(N__13776),
            .I(N__13773));
    LocalMux I__2852 (
            .O(N__13773),
            .I(N__13767));
    CascadeMux I__2851 (
            .O(N__13772),
            .I(N__13763));
    InMux I__2850 (
            .O(N__13771),
            .I(N__13758));
    InMux I__2849 (
            .O(N__13770),
            .I(N__13755));
    Span4Mux_h I__2848 (
            .O(N__13767),
            .I(N__13752));
    InMux I__2847 (
            .O(N__13766),
            .I(N__13749));
    InMux I__2846 (
            .O(N__13763),
            .I(N__13742));
    InMux I__2845 (
            .O(N__13762),
            .I(N__13742));
    InMux I__2844 (
            .O(N__13761),
            .I(N__13742));
    LocalMux I__2843 (
            .O(N__13758),
            .I(\Lab_UT.state_2 ));
    LocalMux I__2842 (
            .O(N__13755),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__2841 (
            .O(N__13752),
            .I(\Lab_UT.state_2 ));
    LocalMux I__2840 (
            .O(N__13749),
            .I(\Lab_UT.state_2 ));
    LocalMux I__2839 (
            .O(N__13742),
            .I(\Lab_UT.state_2 ));
    InMux I__2838 (
            .O(N__13731),
            .I(N__13728));
    LocalMux I__2837 (
            .O(N__13728),
            .I(\Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2 ));
    CascadeMux I__2836 (
            .O(N__13725),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ));
    InMux I__2835 (
            .O(N__13722),
            .I(N__13719));
    LocalMux I__2834 (
            .O(N__13719),
            .I(N__13716));
    Span4Mux_s3_v I__2833 (
            .O(N__13716),
            .I(N__13713));
    Span4Mux_v I__2832 (
            .O(N__13713),
            .I(N__13710));
    Odrv4 I__2831 (
            .O(N__13710),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_1 ));
    InMux I__2830 (
            .O(N__13707),
            .I(N__13704));
    LocalMux I__2829 (
            .O(N__13704),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__2828 (
            .O(N__13701),
            .I(N__13698));
    LocalMux I__2827 (
            .O(N__13698),
            .I(\uu2.m76_am_1 ));
    CascadeMux I__2826 (
            .O(N__13695),
            .I(N__13692));
    InMux I__2825 (
            .O(N__13692),
            .I(N__13689));
    LocalMux I__2824 (
            .O(N__13689),
            .I(\uu2.bitmapZ0Z_84 ));
    InMux I__2823 (
            .O(N__13686),
            .I(N__13683));
    LocalMux I__2822 (
            .O(N__13683),
            .I(N__13680));
    Odrv4 I__2821 (
            .O(N__13680),
            .I(\Lab_UT.bcd2segment1.N_244 ));
    InMux I__2820 (
            .O(N__13677),
            .I(N__13673));
    InMux I__2819 (
            .O(N__13676),
            .I(N__13670));
    LocalMux I__2818 (
            .O(N__13673),
            .I(N__13667));
    LocalMux I__2817 (
            .O(N__13670),
            .I(N__13664));
    Span4Mux_v I__2816 (
            .O(N__13667),
            .I(N__13661));
    Span4Mux_h I__2815 (
            .O(N__13664),
            .I(N__13658));
    Odrv4 I__2814 (
            .O(N__13661),
            .I(\uu2.bitmapZ0Z_168 ));
    Odrv4 I__2813 (
            .O(N__13658),
            .I(\uu2.bitmapZ0Z_168 ));
    CascadeMux I__2812 (
            .O(N__13653),
            .I(\Lab_UT.bcd2segment1.N_246_cascade_ ));
    CascadeMux I__2811 (
            .O(N__13650),
            .I(\Lab_UT.dictrl.un1_state_11_cascade_ ));
    SRMux I__2810 (
            .O(N__13647),
            .I(N__13644));
    LocalMux I__2809 (
            .O(N__13644),
            .I(N__13641));
    Span4Mux_h I__2808 (
            .O(N__13641),
            .I(N__13637));
    InMux I__2807 (
            .O(N__13640),
            .I(N__13634));
    Odrv4 I__2806 (
            .O(N__13637),
            .I(\Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1 ));
    LocalMux I__2805 (
            .O(N__13634),
            .I(\Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1 ));
    InMux I__2804 (
            .O(N__13629),
            .I(N__13623));
    InMux I__2803 (
            .O(N__13628),
            .I(N__13618));
    InMux I__2802 (
            .O(N__13627),
            .I(N__13618));
    InMux I__2801 (
            .O(N__13626),
            .I(N__13615));
    LocalMux I__2800 (
            .O(N__13623),
            .I(N__13612));
    LocalMux I__2799 (
            .O(N__13618),
            .I(N__13609));
    LocalMux I__2798 (
            .O(N__13615),
            .I(N__13602));
    Span4Mux_h I__2797 (
            .O(N__13612),
            .I(N__13602));
    Span4Mux_h I__2796 (
            .O(N__13609),
            .I(N__13602));
    Span4Mux_v I__2795 (
            .O(N__13602),
            .I(N__13599));
    Odrv4 I__2794 (
            .O(N__13599),
            .I(\Lab_UT.bcd2segment1.N_264 ));
    CascadeMux I__2793 (
            .O(N__13596),
            .I(\Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_ ));
    InMux I__2792 (
            .O(N__13593),
            .I(N__13590));
    LocalMux I__2791 (
            .O(N__13590),
            .I(N__13587));
    Span4Mux_h I__2790 (
            .O(N__13587),
            .I(N__13582));
    InMux I__2789 (
            .O(N__13586),
            .I(N__13579));
    InMux I__2788 (
            .O(N__13585),
            .I(N__13576));
    Odrv4 I__2787 (
            .O(N__13582),
            .I(\Lab_UT.dictrl.next_state16Z0Z_5 ));
    LocalMux I__2786 (
            .O(N__13579),
            .I(\Lab_UT.dictrl.next_state16Z0Z_5 ));
    LocalMux I__2785 (
            .O(N__13576),
            .I(\Lab_UT.dictrl.next_state16Z0Z_5 ));
    CascadeMux I__2784 (
            .O(N__13569),
            .I(\Lab_UT.m68_0_ns_cascade_ ));
    InMux I__2783 (
            .O(N__13566),
            .I(N__13561));
    InMux I__2782 (
            .O(N__13565),
            .I(N__13558));
    InMux I__2781 (
            .O(N__13564),
            .I(N__13555));
    LocalMux I__2780 (
            .O(N__13561),
            .I(\Lab_UT.dictrl.next_state16Z0Z_4 ));
    LocalMux I__2779 (
            .O(N__13558),
            .I(\Lab_UT.dictrl.next_state16Z0Z_4 ));
    LocalMux I__2778 (
            .O(N__13555),
            .I(\Lab_UT.dictrl.next_state16Z0Z_4 ));
    InMux I__2777 (
            .O(N__13548),
            .I(N__13545));
    LocalMux I__2776 (
            .O(N__13545),
            .I(N__13539));
    InMux I__2775 (
            .O(N__13544),
            .I(N__13532));
    InMux I__2774 (
            .O(N__13543),
            .I(N__13532));
    InMux I__2773 (
            .O(N__13542),
            .I(N__13532));
    Sp12to4 I__2772 (
            .O(N__13539),
            .I(N__13526));
    LocalMux I__2771 (
            .O(N__13532),
            .I(N__13526));
    InMux I__2770 (
            .O(N__13531),
            .I(N__13523));
    Odrv12 I__2769 (
            .O(N__13526),
            .I(\Lab_UT.state_3 ));
    LocalMux I__2768 (
            .O(N__13523),
            .I(\Lab_UT.state_3 ));
    InMux I__2767 (
            .O(N__13518),
            .I(N__13511));
    InMux I__2766 (
            .O(N__13517),
            .I(N__13511));
    InMux I__2765 (
            .O(N__13516),
            .I(N__13508));
    LocalMux I__2764 (
            .O(N__13511),
            .I(N__13499));
    LocalMux I__2763 (
            .O(N__13508),
            .I(N__13499));
    InMux I__2762 (
            .O(N__13507),
            .I(N__13496));
    InMux I__2761 (
            .O(N__13506),
            .I(N__13489));
    InMux I__2760 (
            .O(N__13505),
            .I(N__13489));
    InMux I__2759 (
            .O(N__13504),
            .I(N__13489));
    Odrv4 I__2758 (
            .O(N__13499),
            .I(\Lab_UT.state_1 ));
    LocalMux I__2757 (
            .O(N__13496),
            .I(\Lab_UT.state_1 ));
    LocalMux I__2756 (
            .O(N__13489),
            .I(\Lab_UT.state_1 ));
    CascadeMux I__2755 (
            .O(N__13482),
            .I(\Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_ ));
    CascadeMux I__2754 (
            .O(N__13479),
            .I(\Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_ ));
    CascadeMux I__2753 (
            .O(N__13476),
            .I(N__13472));
    CascadeMux I__2752 (
            .O(N__13475),
            .I(N__13469));
    InMux I__2751 (
            .O(N__13472),
            .I(N__13466));
    InMux I__2750 (
            .O(N__13469),
            .I(N__13463));
    LocalMux I__2749 (
            .O(N__13466),
            .I(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ));
    LocalMux I__2748 (
            .O(N__13463),
            .I(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ));
    InMux I__2747 (
            .O(N__13458),
            .I(N__13453));
    InMux I__2746 (
            .O(N__13457),
            .I(N__13448));
    InMux I__2745 (
            .O(N__13456),
            .I(N__13448));
    LocalMux I__2744 (
            .O(N__13453),
            .I(N__13445));
    LocalMux I__2743 (
            .O(N__13448),
            .I(N__13442));
    Span4Mux_h I__2742 (
            .O(N__13445),
            .I(N__13439));
    Span4Mux_h I__2741 (
            .O(N__13442),
            .I(N__13436));
    Odrv4 I__2740 (
            .O(N__13439),
            .I(\Lab_UT.dictrl.next_state_set ));
    Odrv4 I__2739 (
            .O(N__13436),
            .I(\Lab_UT.dictrl.next_state_set ));
    CascadeMux I__2738 (
            .O(N__13431),
            .I(\buart.Z_rx.bitcount_lm_3_cascade_ ));
    SRMux I__2737 (
            .O(N__13428),
            .I(N__13424));
    InMux I__2736 (
            .O(N__13427),
            .I(N__13421));
    LocalMux I__2735 (
            .O(N__13424),
            .I(N__13418));
    LocalMux I__2734 (
            .O(N__13421),
            .I(N__13415));
    Odrv12 I__2733 (
            .O(N__13418),
            .I(\Lab_UT.m72_0 ));
    Odrv4 I__2732 (
            .O(N__13415),
            .I(\Lab_UT.m72_0 ));
    InMux I__2731 (
            .O(N__13410),
            .I(N__13400));
    InMux I__2730 (
            .O(N__13409),
            .I(N__13400));
    InMux I__2729 (
            .O(N__13408),
            .I(N__13400));
    InMux I__2728 (
            .O(N__13407),
            .I(N__13397));
    LocalMux I__2727 (
            .O(N__13400),
            .I(N__13394));
    LocalMux I__2726 (
            .O(N__13397),
            .I(\Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1 ));
    Odrv4 I__2725 (
            .O(N__13394),
            .I(\Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1 ));
    CascadeMux I__2724 (
            .O(N__13389),
            .I(N__13386));
    InMux I__2723 (
            .O(N__13386),
            .I(N__13383));
    LocalMux I__2722 (
            .O(N__13383),
            .I(\Lab_UT.un1_state_13 ));
    CascadeMux I__2721 (
            .O(N__13380),
            .I(\Lab_UT.un1_state_13_cascade_ ));
    InMux I__2720 (
            .O(N__13377),
            .I(N__13373));
    InMux I__2719 (
            .O(N__13376),
            .I(N__13370));
    LocalMux I__2718 (
            .O(N__13373),
            .I(N__13365));
    LocalMux I__2717 (
            .O(N__13370),
            .I(N__13365));
    Span4Mux_h I__2716 (
            .O(N__13365),
            .I(N__13362));
    Odrv4 I__2715 (
            .O(N__13362),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__2714 (
            .O(N__13359),
            .I(N__13355));
    InMux I__2713 (
            .O(N__13358),
            .I(N__13352));
    LocalMux I__2712 (
            .O(N__13355),
            .I(N__13349));
    LocalMux I__2711 (
            .O(N__13352),
            .I(N__13346));
    Span4Mux_h I__2710 (
            .O(N__13349),
            .I(N__13343));
    Odrv4 I__2709 (
            .O(N__13346),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__2708 (
            .O(N__13343),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__2707 (
            .O(N__13338),
            .I(N__13335));
    LocalMux I__2706 (
            .O(N__13335),
            .I(\Lab_UT.dictrl.un1_state_11 ));
    CascadeMux I__2705 (
            .O(N__13332),
            .I(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_ ));
    InMux I__2704 (
            .O(N__13329),
            .I(N__13326));
    LocalMux I__2703 (
            .O(N__13326),
            .I(N__13323));
    Span4Mux_v I__2702 (
            .O(N__13323),
            .I(N__13320));
    Odrv4 I__2701 (
            .O(N__13320),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    CascadeMux I__2700 (
            .O(N__13317),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ));
    CascadeMux I__2699 (
            .O(N__13314),
            .I(N__13311));
    InMux I__2698 (
            .O(N__13311),
            .I(N__13308));
    LocalMux I__2697 (
            .O(N__13308),
            .I(N__13305));
    Span4Mux_h I__2696 (
            .O(N__13305),
            .I(N__13301));
    InMux I__2695 (
            .O(N__13304),
            .I(N__13298));
    Odrv4 I__2694 (
            .O(N__13301),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    LocalMux I__2693 (
            .O(N__13298),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    InMux I__2692 (
            .O(N__13293),
            .I(N__13289));
    InMux I__2691 (
            .O(N__13292),
            .I(N__13286));
    LocalMux I__2690 (
            .O(N__13289),
            .I(N__13283));
    LocalMux I__2689 (
            .O(N__13286),
            .I(N__13280));
    Odrv4 I__2688 (
            .O(N__13283),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    Odrv4 I__2687 (
            .O(N__13280),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    CascadeMux I__2686 (
            .O(N__13275),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3_cascade_ ));
    InMux I__2685 (
            .O(N__13272),
            .I(N__13269));
    LocalMux I__2684 (
            .O(N__13269),
            .I(N__13266));
    Span4Mux_h I__2683 (
            .O(N__13266),
            .I(N__13261));
    InMux I__2682 (
            .O(N__13265),
            .I(N__13256));
    InMux I__2681 (
            .O(N__13264),
            .I(N__13256));
    Odrv4 I__2680 (
            .O(N__13261),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    LocalMux I__2679 (
            .O(N__13256),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    InMux I__2678 (
            .O(N__13251),
            .I(N__13248));
    LocalMux I__2677 (
            .O(N__13248),
            .I(N__13245));
    Span4Mux_h I__2676 (
            .O(N__13245),
            .I(N__13242));
    Odrv4 I__2675 (
            .O(N__13242),
            .I(\Lab_UT.dictrl.dicRun_2_reti ));
    InMux I__2674 (
            .O(N__13239),
            .I(N__13236));
    LocalMux I__2673 (
            .O(N__13236),
            .I(\Lab_UT.dictrl.next_state_out_0 ));
    InMux I__2672 (
            .O(N__13233),
            .I(N__13229));
    InMux I__2671 (
            .O(N__13232),
            .I(N__13226));
    LocalMux I__2670 (
            .O(N__13229),
            .I(\uu2.bitmapZ0Z_52 ));
    LocalMux I__2669 (
            .O(N__13226),
            .I(\uu2.bitmapZ0Z_52 ));
    CascadeMux I__2668 (
            .O(N__13221),
            .I(N__13218));
    InMux I__2667 (
            .O(N__13218),
            .I(N__13213));
    InMux I__2666 (
            .O(N__13217),
            .I(N__13210));
    InMux I__2665 (
            .O(N__13216),
            .I(N__13207));
    LocalMux I__2664 (
            .O(N__13213),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__2663 (
            .O(N__13210),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__2662 (
            .O(N__13207),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    CascadeMux I__2661 (
            .O(N__13200),
            .I(\Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_ ));
    CascadeMux I__2660 (
            .O(N__13197),
            .I(\Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_ ));
    InMux I__2659 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__2658 (
            .O(N__13191),
            .I(N__13187));
    CascadeMux I__2657 (
            .O(N__13190),
            .I(N__13184));
    Span4Mux_h I__2656 (
            .O(N__13187),
            .I(N__13179));
    InMux I__2655 (
            .O(N__13184),
            .I(N__13174));
    InMux I__2654 (
            .O(N__13183),
            .I(N__13174));
    InMux I__2653 (
            .O(N__13182),
            .I(N__13171));
    Odrv4 I__2652 (
            .O(N__13179),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    LocalMux I__2651 (
            .O(N__13174),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    LocalMux I__2650 (
            .O(N__13171),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    CascadeMux I__2649 (
            .O(N__13164),
            .I(N__13159));
    InMux I__2648 (
            .O(N__13163),
            .I(N__13155));
    InMux I__2647 (
            .O(N__13162),
            .I(N__13148));
    InMux I__2646 (
            .O(N__13159),
            .I(N__13148));
    InMux I__2645 (
            .O(N__13158),
            .I(N__13148));
    LocalMux I__2644 (
            .O(N__13155),
            .I(N__13145));
    LocalMux I__2643 (
            .O(N__13148),
            .I(N__13142));
    Span4Mux_h I__2642 (
            .O(N__13145),
            .I(N__13139));
    Span4Mux_h I__2641 (
            .O(N__13142),
            .I(N__13136));
    Odrv4 I__2640 (
            .O(N__13139),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv4 I__2639 (
            .O(N__13136),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    CascadeMux I__2638 (
            .O(N__13131),
            .I(N__13127));
    InMux I__2637 (
            .O(N__13130),
            .I(N__13119));
    InMux I__2636 (
            .O(N__13127),
            .I(N__13119));
    InMux I__2635 (
            .O(N__13126),
            .I(N__13119));
    LocalMux I__2634 (
            .O(N__13119),
            .I(N__13116));
    Odrv12 I__2633 (
            .O(N__13116),
            .I(\Lab_UT.N_9_0 ));
    CascadeMux I__2632 (
            .O(N__13113),
            .I(N__13110));
    InMux I__2631 (
            .O(N__13110),
            .I(N__13107));
    LocalMux I__2630 (
            .O(N__13107),
            .I(N__13103));
    CascadeMux I__2629 (
            .O(N__13106),
            .I(N__13099));
    Sp12to4 I__2628 (
            .O(N__13103),
            .I(N__13095));
    InMux I__2627 (
            .O(N__13102),
            .I(N__13088));
    InMux I__2626 (
            .O(N__13099),
            .I(N__13088));
    InMux I__2625 (
            .O(N__13098),
            .I(N__13088));
    Odrv12 I__2624 (
            .O(N__13095),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    LocalMux I__2623 (
            .O(N__13088),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    InMux I__2622 (
            .O(N__13083),
            .I(N__13080));
    LocalMux I__2621 (
            .O(N__13080),
            .I(N__13077));
    Odrv4 I__2620 (
            .O(N__13077),
            .I(\Lab_UT.bcd2segment1.N_181 ));
    InMux I__2619 (
            .O(N__13074),
            .I(N__13071));
    LocalMux I__2618 (
            .O(N__13071),
            .I(N__13068));
    Odrv12 I__2617 (
            .O(N__13068),
            .I(\Lab_UT.bcd2segment1.N_229 ));
    InMux I__2616 (
            .O(N__13065),
            .I(N__13053));
    InMux I__2615 (
            .O(N__13064),
            .I(N__13053));
    InMux I__2614 (
            .O(N__13063),
            .I(N__13053));
    InMux I__2613 (
            .O(N__13062),
            .I(N__13053));
    LocalMux I__2612 (
            .O(N__13053),
            .I(N__13045));
    InMux I__2611 (
            .O(N__13052),
            .I(N__13037));
    InMux I__2610 (
            .O(N__13051),
            .I(N__13037));
    InMux I__2609 (
            .O(N__13050),
            .I(N__13034));
    InMux I__2608 (
            .O(N__13049),
            .I(N__13031));
    InMux I__2607 (
            .O(N__13048),
            .I(N__13028));
    Span4Mux_v I__2606 (
            .O(N__13045),
            .I(N__13025));
    InMux I__2605 (
            .O(N__13044),
            .I(N__13018));
    InMux I__2604 (
            .O(N__13043),
            .I(N__13018));
    InMux I__2603 (
            .O(N__13042),
            .I(N__13018));
    LocalMux I__2602 (
            .O(N__13037),
            .I(N__13015));
    LocalMux I__2601 (
            .O(N__13034),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__2600 (
            .O(N__13031),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__2599 (
            .O(N__13028),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__2598 (
            .O(N__13025),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__2597 (
            .O(N__13018),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__2596 (
            .O(N__13015),
            .I(\Lab_UT.di_Mtens_3 ));
    InMux I__2595 (
            .O(N__13002),
            .I(N__12990));
    InMux I__2594 (
            .O(N__13001),
            .I(N__12990));
    InMux I__2593 (
            .O(N__13000),
            .I(N__12990));
    InMux I__2592 (
            .O(N__12999),
            .I(N__12990));
    LocalMux I__2591 (
            .O(N__12990),
            .I(N__12982));
    InMux I__2590 (
            .O(N__12989),
            .I(N__12973));
    InMux I__2589 (
            .O(N__12988),
            .I(N__12973));
    InMux I__2588 (
            .O(N__12987),
            .I(N__12973));
    InMux I__2587 (
            .O(N__12986),
            .I(N__12973));
    InMux I__2586 (
            .O(N__12985),
            .I(N__12968));
    Span4Mux_h I__2585 (
            .O(N__12982),
            .I(N__12963));
    LocalMux I__2584 (
            .O(N__12973),
            .I(N__12960));
    InMux I__2583 (
            .O(N__12972),
            .I(N__12954));
    InMux I__2582 (
            .O(N__12971),
            .I(N__12954));
    LocalMux I__2581 (
            .O(N__12968),
            .I(N__12951));
    InMux I__2580 (
            .O(N__12967),
            .I(N__12946));
    InMux I__2579 (
            .O(N__12966),
            .I(N__12946));
    Sp12to4 I__2578 (
            .O(N__12963),
            .I(N__12943));
    Span4Mux_h I__2577 (
            .O(N__12960),
            .I(N__12940));
    InMux I__2576 (
            .O(N__12959),
            .I(N__12937));
    LocalMux I__2575 (
            .O(N__12954),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__2574 (
            .O(N__12951),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__2573 (
            .O(N__12946),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv12 I__2572 (
            .O(N__12943),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__2571 (
            .O(N__12940),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__2570 (
            .O(N__12937),
            .I(\Lab_UT.di_Mtens_1 ));
    CascadeMux I__2569 (
            .O(N__12924),
            .I(N__12917));
    InMux I__2568 (
            .O(N__12923),
            .I(N__12914));
    InMux I__2567 (
            .O(N__12922),
            .I(N__12903));
    InMux I__2566 (
            .O(N__12921),
            .I(N__12903));
    InMux I__2565 (
            .O(N__12920),
            .I(N__12903));
    InMux I__2564 (
            .O(N__12917),
            .I(N__12903));
    LocalMux I__2563 (
            .O(N__12914),
            .I(N__12898));
    InMux I__2562 (
            .O(N__12913),
            .I(N__12893));
    InMux I__2561 (
            .O(N__12912),
            .I(N__12893));
    LocalMux I__2560 (
            .O(N__12903),
            .I(N__12890));
    CascadeMux I__2559 (
            .O(N__12902),
            .I(N__12884));
    CascadeMux I__2558 (
            .O(N__12901),
            .I(N__12880));
    Span4Mux_h I__2557 (
            .O(N__12898),
            .I(N__12877));
    LocalMux I__2556 (
            .O(N__12893),
            .I(N__12872));
    Span12Mux_s9_v I__2555 (
            .O(N__12890),
            .I(N__12872));
    InMux I__2554 (
            .O(N__12889),
            .I(N__12863));
    InMux I__2553 (
            .O(N__12888),
            .I(N__12863));
    InMux I__2552 (
            .O(N__12887),
            .I(N__12863));
    InMux I__2551 (
            .O(N__12884),
            .I(N__12863));
    InMux I__2550 (
            .O(N__12883),
            .I(N__12858));
    InMux I__2549 (
            .O(N__12880),
            .I(N__12858));
    Odrv4 I__2548 (
            .O(N__12877),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv12 I__2547 (
            .O(N__12872),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__2546 (
            .O(N__12863),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__2545 (
            .O(N__12858),
            .I(\Lab_UT.di_Mtens_2 ));
    InMux I__2544 (
            .O(N__12849),
            .I(N__12846));
    LocalMux I__2543 (
            .O(N__12846),
            .I(N__12843));
    Odrv4 I__2542 (
            .O(N__12843),
            .I(\Lab_UT.bcd2segment1.N_233 ));
    InMux I__2541 (
            .O(N__12840),
            .I(N__12836));
    InMux I__2540 (
            .O(N__12839),
            .I(N__12833));
    LocalMux I__2539 (
            .O(N__12836),
            .I(N__12829));
    LocalMux I__2538 (
            .O(N__12833),
            .I(N__12826));
    InMux I__2537 (
            .O(N__12832),
            .I(N__12823));
    Span4Mux_h I__2536 (
            .O(N__12829),
            .I(N__12820));
    Span4Mux_h I__2535 (
            .O(N__12826),
            .I(N__12817));
    LocalMux I__2534 (
            .O(N__12823),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__2533 (
            .O(N__12820),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__2532 (
            .O(N__12817),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    CascadeMux I__2531 (
            .O(N__12810),
            .I(N__12804));
    InMux I__2530 (
            .O(N__12809),
            .I(N__12797));
    InMux I__2529 (
            .O(N__12808),
            .I(N__12797));
    InMux I__2528 (
            .O(N__12807),
            .I(N__12797));
    InMux I__2527 (
            .O(N__12804),
            .I(N__12794));
    LocalMux I__2526 (
            .O(N__12797),
            .I(N__12791));
    LocalMux I__2525 (
            .O(N__12794),
            .I(N__12788));
    Span4Mux_h I__2524 (
            .O(N__12791),
            .I(N__12785));
    Span4Mux_h I__2523 (
            .O(N__12788),
            .I(N__12782));
    Odrv4 I__2522 (
            .O(N__12785),
            .I(\uu2.N_115 ));
    Odrv4 I__2521 (
            .O(N__12782),
            .I(\uu2.N_115 ));
    CascadeMux I__2520 (
            .O(N__12777),
            .I(N__12773));
    InMux I__2519 (
            .O(N__12776),
            .I(N__12763));
    InMux I__2518 (
            .O(N__12773),
            .I(N__12763));
    InMux I__2517 (
            .O(N__12772),
            .I(N__12763));
    CascadeMux I__2516 (
            .O(N__12771),
            .I(N__12760));
    CascadeMux I__2515 (
            .O(N__12770),
            .I(N__12756));
    LocalMux I__2514 (
            .O(N__12763),
            .I(N__12750));
    InMux I__2513 (
            .O(N__12760),
            .I(N__12747));
    InMux I__2512 (
            .O(N__12759),
            .I(N__12744));
    InMux I__2511 (
            .O(N__12756),
            .I(N__12741));
    CascadeMux I__2510 (
            .O(N__12755),
            .I(N__12738));
    CascadeMux I__2509 (
            .O(N__12754),
            .I(N__12733));
    CascadeMux I__2508 (
            .O(N__12753),
            .I(N__12728));
    Span4Mux_v I__2507 (
            .O(N__12750),
            .I(N__12722));
    LocalMux I__2506 (
            .O(N__12747),
            .I(N__12722));
    LocalMux I__2505 (
            .O(N__12744),
            .I(N__12717));
    LocalMux I__2504 (
            .O(N__12741),
            .I(N__12717));
    InMux I__2503 (
            .O(N__12738),
            .I(N__12710));
    InMux I__2502 (
            .O(N__12737),
            .I(N__12710));
    InMux I__2501 (
            .O(N__12736),
            .I(N__12710));
    InMux I__2500 (
            .O(N__12733),
            .I(N__12707));
    InMux I__2499 (
            .O(N__12732),
            .I(N__12700));
    InMux I__2498 (
            .O(N__12731),
            .I(N__12700));
    InMux I__2497 (
            .O(N__12728),
            .I(N__12700));
    InMux I__2496 (
            .O(N__12727),
            .I(N__12697));
    Span4Mux_h I__2495 (
            .O(N__12722),
            .I(N__12694));
    Span4Mux_h I__2494 (
            .O(N__12717),
            .I(N__12691));
    LocalMux I__2493 (
            .O(N__12710),
            .I(N__12686));
    LocalMux I__2492 (
            .O(N__12707),
            .I(N__12686));
    LocalMux I__2491 (
            .O(N__12700),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2490 (
            .O(N__12697),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2489 (
            .O(N__12694),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2488 (
            .O(N__12691),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2487 (
            .O(N__12686),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    CascadeMux I__2486 (
            .O(N__12675),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_ ));
    InMux I__2485 (
            .O(N__12672),
            .I(N__12669));
    LocalMux I__2484 (
            .O(N__12669),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_0 ));
    CascadeMux I__2483 (
            .O(N__12666),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_ ));
    CascadeMux I__2482 (
            .O(N__12663),
            .I(N__12660));
    InMux I__2481 (
            .O(N__12660),
            .I(N__12657));
    LocalMux I__2480 (
            .O(N__12657),
            .I(N__12654));
    Odrv12 I__2479 (
            .O(N__12654),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__2478 (
            .O(N__12651),
            .I(N__12647));
    InMux I__2477 (
            .O(N__12650),
            .I(N__12644));
    LocalMux I__2476 (
            .O(N__12647),
            .I(\uu2.bitmapZ0Z_308 ));
    LocalMux I__2475 (
            .O(N__12644),
            .I(\uu2.bitmapZ0Z_308 ));
    CascadeMux I__2474 (
            .O(N__12639),
            .I(\uu2.mem0.m317_0_a6_0_cascade_ ));
    InMux I__2473 (
            .O(N__12636),
            .I(N__12633));
    LocalMux I__2472 (
            .O(N__12633),
            .I(N__12630));
    Odrv4 I__2471 (
            .O(N__12630),
            .I(\uu2.mem0.N_6_0 ));
    InMux I__2470 (
            .O(N__12627),
            .I(N__12624));
    LocalMux I__2469 (
            .O(N__12624),
            .I(\uu2.mem0.m317_0_0 ));
    CascadeMux I__2468 (
            .O(N__12621),
            .I(\uu2.mem0.N_11_0_0_cascade_ ));
    InMux I__2467 (
            .O(N__12618),
            .I(N__12615));
    LocalMux I__2466 (
            .O(N__12615),
            .I(N__12612));
    Odrv4 I__2465 (
            .O(N__12612),
            .I(\uu2.mem0.N_6_0_0_0 ));
    InMux I__2464 (
            .O(N__12609),
            .I(N__12602));
    InMux I__2463 (
            .O(N__12608),
            .I(N__12602));
    CascadeMux I__2462 (
            .O(N__12607),
            .I(N__12596));
    LocalMux I__2461 (
            .O(N__12602),
            .I(N__12591));
    InMux I__2460 (
            .O(N__12601),
            .I(N__12582));
    InMux I__2459 (
            .O(N__12600),
            .I(N__12582));
    InMux I__2458 (
            .O(N__12599),
            .I(N__12582));
    InMux I__2457 (
            .O(N__12596),
            .I(N__12582));
    InMux I__2456 (
            .O(N__12595),
            .I(N__12577));
    InMux I__2455 (
            .O(N__12594),
            .I(N__12577));
    Odrv4 I__2454 (
            .O(N__12591),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__2453 (
            .O(N__12582),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__2452 (
            .O(N__12577),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    InMux I__2451 (
            .O(N__12570),
            .I(N__12567));
    LocalMux I__2450 (
            .O(N__12567),
            .I(\uu2.mem0.N_5_0 ));
    InMux I__2449 (
            .O(N__12564),
            .I(N__12561));
    LocalMux I__2448 (
            .O(N__12561),
            .I(\uu2.mem0.N_14 ));
    InMux I__2447 (
            .O(N__12558),
            .I(N__12555));
    LocalMux I__2446 (
            .O(N__12555),
            .I(N__12552));
    Odrv12 I__2445 (
            .O(N__12552),
            .I(\uu2.mem0.g1_2_2_2_1 ));
    InMux I__2444 (
            .O(N__12549),
            .I(N__12545));
    InMux I__2443 (
            .O(N__12548),
            .I(N__12542));
    LocalMux I__2442 (
            .O(N__12545),
            .I(\uu2.bitmapZ0Z_34 ));
    LocalMux I__2441 (
            .O(N__12542),
            .I(\uu2.bitmapZ0Z_34 ));
    InMux I__2440 (
            .O(N__12537),
            .I(N__12534));
    LocalMux I__2439 (
            .O(N__12534),
            .I(N__12531));
    Span4Mux_v I__2438 (
            .O(N__12531),
            .I(N__12528));
    Odrv4 I__2437 (
            .O(N__12528),
            .I(\Lab_UT.bcd2segment1.N_239 ));
    InMux I__2436 (
            .O(N__12525),
            .I(N__12521));
    InMux I__2435 (
            .O(N__12524),
            .I(N__12518));
    LocalMux I__2434 (
            .O(N__12521),
            .I(\uu2.bitmapZ0Z_290 ));
    LocalMux I__2433 (
            .O(N__12518),
            .I(\uu2.bitmapZ0Z_290 ));
    CascadeMux I__2432 (
            .O(N__12513),
            .I(N__12508));
    InMux I__2431 (
            .O(N__12512),
            .I(N__12505));
    InMux I__2430 (
            .O(N__12511),
            .I(N__12500));
    InMux I__2429 (
            .O(N__12508),
            .I(N__12500));
    LocalMux I__2428 (
            .O(N__12505),
            .I(N__12495));
    LocalMux I__2427 (
            .O(N__12500),
            .I(N__12495));
    Odrv12 I__2426 (
            .O(N__12495),
            .I(\uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8 ));
    InMux I__2425 (
            .O(N__12492),
            .I(N__12488));
    InMux I__2424 (
            .O(N__12491),
            .I(N__12485));
    LocalMux I__2423 (
            .O(N__12488),
            .I(N__12482));
    LocalMux I__2422 (
            .O(N__12485),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    Odrv4 I__2421 (
            .O(N__12482),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    CascadeMux I__2420 (
            .O(N__12477),
            .I(N__12468));
    InMux I__2419 (
            .O(N__12476),
            .I(N__12465));
    InMux I__2418 (
            .O(N__12475),
            .I(N__12462));
    InMux I__2417 (
            .O(N__12474),
            .I(N__12459));
    InMux I__2416 (
            .O(N__12473),
            .I(N__12456));
    InMux I__2415 (
            .O(N__12472),
            .I(N__12453));
    InMux I__2414 (
            .O(N__12471),
            .I(N__12448));
    InMux I__2413 (
            .O(N__12468),
            .I(N__12448));
    LocalMux I__2412 (
            .O(N__12465),
            .I(N__12444));
    LocalMux I__2411 (
            .O(N__12462),
            .I(N__12441));
    LocalMux I__2410 (
            .O(N__12459),
            .I(N__12434));
    LocalMux I__2409 (
            .O(N__12456),
            .I(N__12434));
    LocalMux I__2408 (
            .O(N__12453),
            .I(N__12434));
    LocalMux I__2407 (
            .O(N__12448),
            .I(N__12429));
    InMux I__2406 (
            .O(N__12447),
            .I(N__12421));
    Span4Mux_h I__2405 (
            .O(N__12444),
            .I(N__12418));
    Span4Mux_h I__2404 (
            .O(N__12441),
            .I(N__12415));
    Span4Mux_v I__2403 (
            .O(N__12434),
            .I(N__12412));
    InMux I__2402 (
            .O(N__12433),
            .I(N__12409));
    InMux I__2401 (
            .O(N__12432),
            .I(N__12406));
    Span4Mux_h I__2400 (
            .O(N__12429),
            .I(N__12403));
    InMux I__2399 (
            .O(N__12428),
            .I(N__12398));
    InMux I__2398 (
            .O(N__12427),
            .I(N__12398));
    InMux I__2397 (
            .O(N__12426),
            .I(N__12391));
    InMux I__2396 (
            .O(N__12425),
            .I(N__12391));
    InMux I__2395 (
            .O(N__12424),
            .I(N__12391));
    LocalMux I__2394 (
            .O(N__12421),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2393 (
            .O(N__12418),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2392 (
            .O(N__12415),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2391 (
            .O(N__12412),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2390 (
            .O(N__12409),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2389 (
            .O(N__12406),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2388 (
            .O(N__12403),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2387 (
            .O(N__12398),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2386 (
            .O(N__12391),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    InMux I__2385 (
            .O(N__12372),
            .I(N__12369));
    LocalMux I__2384 (
            .O(N__12369),
            .I(N__12364));
    InMux I__2383 (
            .O(N__12368),
            .I(N__12361));
    CascadeMux I__2382 (
            .O(N__12367),
            .I(N__12355));
    Span4Mux_h I__2381 (
            .O(N__12364),
            .I(N__12348));
    LocalMux I__2380 (
            .O(N__12361),
            .I(N__12348));
    InMux I__2379 (
            .O(N__12360),
            .I(N__12345));
    InMux I__2378 (
            .O(N__12359),
            .I(N__12342));
    InMux I__2377 (
            .O(N__12358),
            .I(N__12332));
    InMux I__2376 (
            .O(N__12355),
            .I(N__12332));
    InMux I__2375 (
            .O(N__12354),
            .I(N__12332));
    InMux I__2374 (
            .O(N__12353),
            .I(N__12332));
    Span4Mux_h I__2373 (
            .O(N__12348),
            .I(N__12321));
    LocalMux I__2372 (
            .O(N__12345),
            .I(N__12316));
    LocalMux I__2371 (
            .O(N__12342),
            .I(N__12316));
    InMux I__2370 (
            .O(N__12341),
            .I(N__12313));
    LocalMux I__2369 (
            .O(N__12332),
            .I(N__12310));
    InMux I__2368 (
            .O(N__12331),
            .I(N__12303));
    InMux I__2367 (
            .O(N__12330),
            .I(N__12303));
    InMux I__2366 (
            .O(N__12329),
            .I(N__12303));
    InMux I__2365 (
            .O(N__12328),
            .I(N__12300));
    InMux I__2364 (
            .O(N__12327),
            .I(N__12293));
    InMux I__2363 (
            .O(N__12326),
            .I(N__12293));
    InMux I__2362 (
            .O(N__12325),
            .I(N__12293));
    InMux I__2361 (
            .O(N__12324),
            .I(N__12290));
    Span4Mux_v I__2360 (
            .O(N__12321),
            .I(N__12287));
    Span4Mux_h I__2359 (
            .O(N__12316),
            .I(N__12282));
    LocalMux I__2358 (
            .O(N__12313),
            .I(N__12282));
    Span4Mux_h I__2357 (
            .O(N__12310),
            .I(N__12279));
    LocalMux I__2356 (
            .O(N__12303),
            .I(N__12276));
    LocalMux I__2355 (
            .O(N__12300),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2354 (
            .O(N__12293),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2353 (
            .O(N__12290),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2352 (
            .O(N__12287),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2351 (
            .O(N__12282),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2350 (
            .O(N__12279),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2349 (
            .O(N__12276),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__2348 (
            .O(N__12261),
            .I(N__12258));
    LocalMux I__2347 (
            .O(N__12258),
            .I(N__12254));
    InMux I__2346 (
            .O(N__12257),
            .I(N__12251));
    Odrv12 I__2345 (
            .O(N__12254),
            .I(\uu2.N_9_i ));
    LocalMux I__2344 (
            .O(N__12251),
            .I(\uu2.N_9_i ));
    InMux I__2343 (
            .O(N__12246),
            .I(N__12242));
    InMux I__2342 (
            .O(N__12245),
            .I(N__12239));
    LocalMux I__2341 (
            .O(N__12242),
            .I(N__12234));
    LocalMux I__2340 (
            .O(N__12239),
            .I(N__12234));
    Odrv12 I__2339 (
            .O(N__12234),
            .I(\uu2.bitmapZ0Z_162 ));
    CascadeMux I__2338 (
            .O(N__12231),
            .I(\uu2.mem0.N_9_cascade_ ));
    InMux I__2337 (
            .O(N__12228),
            .I(N__12225));
    LocalMux I__2336 (
            .O(N__12225),
            .I(\uu2.mem0.N_15 ));
    InMux I__2335 (
            .O(N__12222),
            .I(N__12217));
    CascadeMux I__2334 (
            .O(N__12221),
            .I(N__12210));
    InMux I__2333 (
            .O(N__12220),
            .I(N__12204));
    LocalMux I__2332 (
            .O(N__12217),
            .I(N__12201));
    InMux I__2331 (
            .O(N__12216),
            .I(N__12196));
    InMux I__2330 (
            .O(N__12215),
            .I(N__12196));
    InMux I__2329 (
            .O(N__12214),
            .I(N__12193));
    InMux I__2328 (
            .O(N__12213),
            .I(N__12188));
    InMux I__2327 (
            .O(N__12210),
            .I(N__12188));
    InMux I__2326 (
            .O(N__12209),
            .I(N__12181));
    InMux I__2325 (
            .O(N__12208),
            .I(N__12181));
    InMux I__2324 (
            .O(N__12207),
            .I(N__12181));
    LocalMux I__2323 (
            .O(N__12204),
            .I(N__12178));
    Span4Mux_v I__2322 (
            .O(N__12201),
            .I(N__12173));
    LocalMux I__2321 (
            .O(N__12196),
            .I(N__12173));
    LocalMux I__2320 (
            .O(N__12193),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2319 (
            .O(N__12188),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2318 (
            .O(N__12181),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv12 I__2317 (
            .O(N__12178),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__2316 (
            .O(N__12173),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__2315 (
            .O(N__12162),
            .I(N__12159));
    LocalMux I__2314 (
            .O(N__12159),
            .I(N__12156));
    Odrv4 I__2313 (
            .O(N__12156),
            .I(\uu2.mem0.N_7 ));
    CascadeMux I__2312 (
            .O(N__12153),
            .I(\uu2.N_126_cascade_ ));
    InMux I__2311 (
            .O(N__12150),
            .I(N__12143));
    InMux I__2310 (
            .O(N__12149),
            .I(N__12139));
    InMux I__2309 (
            .O(N__12148),
            .I(N__12136));
    InMux I__2308 (
            .O(N__12147),
            .I(N__12131));
    InMux I__2307 (
            .O(N__12146),
            .I(N__12131));
    LocalMux I__2306 (
            .O(N__12143),
            .I(N__12128));
    InMux I__2305 (
            .O(N__12142),
            .I(N__12125));
    LocalMux I__2304 (
            .O(N__12139),
            .I(N__12120));
    LocalMux I__2303 (
            .O(N__12136),
            .I(N__12120));
    LocalMux I__2302 (
            .O(N__12131),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv12 I__2301 (
            .O(N__12128),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__2300 (
            .O(N__12125),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__2299 (
            .O(N__12120),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__2298 (
            .O(N__12111),
            .I(N__12108));
    InMux I__2297 (
            .O(N__12108),
            .I(N__12105));
    LocalMux I__2296 (
            .O(N__12105),
            .I(N__12102));
    Odrv12 I__2295 (
            .O(N__12102),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0 ));
    InMux I__2294 (
            .O(N__12099),
            .I(N__12096));
    LocalMux I__2293 (
            .O(N__12096),
            .I(N__12093));
    Span4Mux_v I__2292 (
            .O(N__12093),
            .I(N__12090));
    Odrv4 I__2291 (
            .O(N__12090),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_67 ));
    InMux I__2290 (
            .O(N__12087),
            .I(N__12084));
    LocalMux I__2289 (
            .O(N__12084),
            .I(N__12081));
    Span4Mux_h I__2288 (
            .O(N__12081),
            .I(N__12078));
    Odrv4 I__2287 (
            .O(N__12078),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_66 ));
    InMux I__2286 (
            .O(N__12075),
            .I(N__12071));
    InMux I__2285 (
            .O(N__12074),
            .I(N__12068));
    LocalMux I__2284 (
            .O(N__12071),
            .I(N__12065));
    LocalMux I__2283 (
            .O(N__12068),
            .I(N__12060));
    Span4Mux_h I__2282 (
            .O(N__12065),
            .I(N__12057));
    InMux I__2281 (
            .O(N__12064),
            .I(N__12052));
    InMux I__2280 (
            .O(N__12063),
            .I(N__12052));
    Odrv12 I__2279 (
            .O(N__12060),
            .I(\uu2.N_126 ));
    Odrv4 I__2278 (
            .O(N__12057),
            .I(\uu2.N_126 ));
    LocalMux I__2277 (
            .O(N__12052),
            .I(\uu2.N_126 ));
    InMux I__2276 (
            .O(N__12045),
            .I(N__12042));
    LocalMux I__2275 (
            .O(N__12042),
            .I(N__12039));
    Span4Mux_v I__2274 (
            .O(N__12039),
            .I(N__12036));
    Span4Mux_h I__2273 (
            .O(N__12036),
            .I(N__12033));
    Odrv4 I__2272 (
            .O(N__12033),
            .I(\uu2.mem0.g0_7_0_0 ));
    CascadeMux I__2271 (
            .O(N__12030),
            .I(\uu2.mem0.N_57_cascade_ ));
    InMux I__2270 (
            .O(N__12027),
            .I(N__12024));
    LocalMux I__2269 (
            .O(N__12024),
            .I(\uu2.mem0.bitmap_pmux_u_i_5_1 ));
    InMux I__2268 (
            .O(N__12021),
            .I(N__12018));
    LocalMux I__2267 (
            .O(N__12018),
            .I(\uu2.mem0.g0_7_0_3 ));
    InMux I__2266 (
            .O(N__12015),
            .I(N__12012));
    LocalMux I__2265 (
            .O(N__12012),
            .I(\uu2.N_16 ));
    CascadeMux I__2264 (
            .O(N__12009),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_ ));
    InMux I__2263 (
            .O(N__12006),
            .I(N__12003));
    LocalMux I__2262 (
            .O(N__12003),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_57 ));
    InMux I__2261 (
            .O(N__12000),
            .I(N__11997));
    LocalMux I__2260 (
            .O(N__11997),
            .I(\uu2.mem0.N_13_0 ));
    InMux I__2259 (
            .O(N__11994),
            .I(N__11990));
    InMux I__2258 (
            .O(N__11993),
            .I(N__11987));
    LocalMux I__2257 (
            .O(N__11990),
            .I(\uu2.N_8 ));
    LocalMux I__2256 (
            .O(N__11987),
            .I(\uu2.N_8 ));
    CascadeMux I__2255 (
            .O(N__11982),
            .I(\Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_ ));
    CascadeMux I__2254 (
            .O(N__11979),
            .I(\uu2.N_1580_0_cascade_ ));
    InMux I__2253 (
            .O(N__11976),
            .I(N__11973));
    LocalMux I__2252 (
            .O(N__11973),
            .I(N__11969));
    CascadeMux I__2251 (
            .O(N__11972),
            .I(N__11966));
    Span4Mux_h I__2250 (
            .O(N__11969),
            .I(N__11963));
    InMux I__2249 (
            .O(N__11966),
            .I(N__11960));
    Odrv4 I__2248 (
            .O(N__11963),
            .I(\uu2.N_77_0 ));
    LocalMux I__2247 (
            .O(N__11960),
            .I(\uu2.N_77_0 ));
    InMux I__2246 (
            .O(N__11955),
            .I(N__11947));
    InMux I__2245 (
            .O(N__11954),
            .I(N__11947));
    InMux I__2244 (
            .O(N__11953),
            .I(N__11944));
    InMux I__2243 (
            .O(N__11952),
            .I(N__11940));
    LocalMux I__2242 (
            .O(N__11947),
            .I(N__11933));
    LocalMux I__2241 (
            .O(N__11944),
            .I(N__11930));
    InMux I__2240 (
            .O(N__11943),
            .I(N__11927));
    LocalMux I__2239 (
            .O(N__11940),
            .I(N__11924));
    InMux I__2238 (
            .O(N__11939),
            .I(N__11919));
    InMux I__2237 (
            .O(N__11938),
            .I(N__11919));
    InMux I__2236 (
            .O(N__11937),
            .I(N__11914));
    InMux I__2235 (
            .O(N__11936),
            .I(N__11914));
    Span4Mux_h I__2234 (
            .O(N__11933),
            .I(N__11911));
    Span4Mux_h I__2233 (
            .O(N__11930),
            .I(N__11908));
    LocalMux I__2232 (
            .O(N__11927),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__2231 (
            .O(N__11924),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__2230 (
            .O(N__11919),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__2229 (
            .O(N__11914),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__2228 (
            .O(N__11911),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__2227 (
            .O(N__11908),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__2226 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__2225 (
            .O(N__11892),
            .I(\uu2.bitmapZ0Z_75 ));
    CascadeMux I__2224 (
            .O(N__11889),
            .I(N__11886));
    InMux I__2223 (
            .O(N__11886),
            .I(N__11883));
    LocalMux I__2222 (
            .O(N__11883),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__2221 (
            .O(N__11880),
            .I(N__11877));
    LocalMux I__2220 (
            .O(N__11877),
            .I(\uu2.N_1581_0 ));
    InMux I__2219 (
            .O(N__11874),
            .I(N__11871));
    LocalMux I__2218 (
            .O(N__11871),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__2217 (
            .O(N__11868),
            .I(N__11865));
    LocalMux I__2216 (
            .O(N__11865),
            .I(N__11862));
    Span4Mux_h I__2215 (
            .O(N__11862),
            .I(N__11857));
    InMux I__2214 (
            .O(N__11861),
            .I(N__11852));
    InMux I__2213 (
            .O(N__11860),
            .I(N__11852));
    Odrv4 I__2212 (
            .O(N__11857),
            .I(L3_tx_data_5));
    LocalMux I__2211 (
            .O(N__11852),
            .I(L3_tx_data_5));
    CascadeMux I__2210 (
            .O(N__11847),
            .I(\uu2.mem0.N_134_mux_cascade_ ));
    InMux I__2209 (
            .O(N__11844),
            .I(N__11840));
    InMux I__2208 (
            .O(N__11843),
            .I(N__11837));
    LocalMux I__2207 (
            .O(N__11840),
            .I(N__11831));
    LocalMux I__2206 (
            .O(N__11837),
            .I(N__11828));
    InMux I__2205 (
            .O(N__11836),
            .I(N__11821));
    InMux I__2204 (
            .O(N__11835),
            .I(N__11821));
    InMux I__2203 (
            .O(N__11834),
            .I(N__11821));
    Span4Mux_h I__2202 (
            .O(N__11831),
            .I(N__11818));
    Span4Mux_h I__2201 (
            .O(N__11828),
            .I(N__11813));
    LocalMux I__2200 (
            .O(N__11821),
            .I(N__11813));
    Odrv4 I__2199 (
            .O(N__11818),
            .I(\uu2.w_data_i_0_tzZ0Z_0 ));
    Odrv4 I__2198 (
            .O(N__11813),
            .I(\uu2.w_data_i_0_tzZ0Z_0 ));
    InMux I__2197 (
            .O(N__11808),
            .I(N__11805));
    LocalMux I__2196 (
            .O(N__11805),
            .I(N__11802));
    Span12Mux_s7_h I__2195 (
            .O(N__11802),
            .I(N__11799));
    Odrv12 I__2194 (
            .O(N__11799),
            .I(\uu2.mem0.N_60_0_i ));
    InMux I__2193 (
            .O(N__11796),
            .I(N__11793));
    LocalMux I__2192 (
            .O(N__11793),
            .I(\uu2.mem0.N_55_0 ));
    CascadeMux I__2191 (
            .O(N__11790),
            .I(\Lab_UT.bcd2segment1.N_127_mux_cascade_ ));
    CascadeMux I__2190 (
            .O(N__11787),
            .I(\Lab_UT.bcd2segment1.N_235_cascade_ ));
    CascadeMux I__2189 (
            .O(N__11784),
            .I(\Lab_UT.bcd2segment1.N_237_cascade_ ));
    InMux I__2188 (
            .O(N__11781),
            .I(N__11778));
    LocalMux I__2187 (
            .O(N__11778),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__2186 (
            .O(N__11775),
            .I(N__11772));
    LocalMux I__2185 (
            .O(N__11772),
            .I(\uu2.bitmapZ0Z_194 ));
    InMux I__2184 (
            .O(N__11769),
            .I(N__11763));
    InMux I__2183 (
            .O(N__11768),
            .I(N__11763));
    LocalMux I__2182 (
            .O(N__11763),
            .I(\uu2.N_101_0 ));
    CascadeMux I__2181 (
            .O(N__11760),
            .I(\Lab_UT.bcd2segment1.N_242_cascade_ ));
    InMux I__2180 (
            .O(N__11757),
            .I(N__11754));
    LocalMux I__2179 (
            .O(N__11754),
            .I(N__11751));
    Odrv12 I__2178 (
            .O(N__11751),
            .I(\resetGen.escKeyZ0Z_5 ));
    InMux I__2177 (
            .O(N__11748),
            .I(N__11745));
    LocalMux I__2176 (
            .O(N__11745),
            .I(\Lab_UT.dictrl.next_state_set_0_1 ));
    CascadeMux I__2175 (
            .O(N__11742),
            .I(N__11737));
    InMux I__2174 (
            .O(N__11741),
            .I(N__11734));
    InMux I__2173 (
            .O(N__11740),
            .I(N__11728));
    InMux I__2172 (
            .O(N__11737),
            .I(N__11725));
    LocalMux I__2171 (
            .O(N__11734),
            .I(N__11722));
    InMux I__2170 (
            .O(N__11733),
            .I(N__11715));
    InMux I__2169 (
            .O(N__11732),
            .I(N__11715));
    InMux I__2168 (
            .O(N__11731),
            .I(N__11715));
    LocalMux I__2167 (
            .O(N__11728),
            .I(bu_rx_data_6));
    LocalMux I__2166 (
            .O(N__11725),
            .I(bu_rx_data_6));
    Odrv4 I__2165 (
            .O(N__11722),
            .I(bu_rx_data_6));
    LocalMux I__2164 (
            .O(N__11715),
            .I(bu_rx_data_6));
    CascadeMux I__2163 (
            .O(N__11706),
            .I(N__11699));
    CascadeMux I__2162 (
            .O(N__11705),
            .I(N__11696));
    CascadeMux I__2161 (
            .O(N__11704),
            .I(N__11693));
    CascadeMux I__2160 (
            .O(N__11703),
            .I(N__11689));
    InMux I__2159 (
            .O(N__11702),
            .I(N__11684));
    InMux I__2158 (
            .O(N__11699),
            .I(N__11684));
    InMux I__2157 (
            .O(N__11696),
            .I(N__11681));
    InMux I__2156 (
            .O(N__11693),
            .I(N__11674));
    InMux I__2155 (
            .O(N__11692),
            .I(N__11674));
    InMux I__2154 (
            .O(N__11689),
            .I(N__11674));
    LocalMux I__2153 (
            .O(N__11684),
            .I(bu_rx_data_7));
    LocalMux I__2152 (
            .O(N__11681),
            .I(bu_rx_data_7));
    LocalMux I__2151 (
            .O(N__11674),
            .I(bu_rx_data_7));
    InMux I__2150 (
            .O(N__11667),
            .I(N__11662));
    CascadeMux I__2149 (
            .O(N__11666),
            .I(N__11657));
    InMux I__2148 (
            .O(N__11665),
            .I(N__11653));
    LocalMux I__2147 (
            .O(N__11662),
            .I(N__11650));
    InMux I__2146 (
            .O(N__11661),
            .I(N__11647));
    InMux I__2145 (
            .O(N__11660),
            .I(N__11640));
    InMux I__2144 (
            .O(N__11657),
            .I(N__11640));
    InMux I__2143 (
            .O(N__11656),
            .I(N__11640));
    LocalMux I__2142 (
            .O(N__11653),
            .I(bu_rx_data_4));
    Odrv4 I__2141 (
            .O(N__11650),
            .I(bu_rx_data_4));
    LocalMux I__2140 (
            .O(N__11647),
            .I(bu_rx_data_4));
    LocalMux I__2139 (
            .O(N__11640),
            .I(bu_rx_data_4));
    InMux I__2138 (
            .O(N__11631),
            .I(N__11628));
    LocalMux I__2137 (
            .O(N__11628),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0 ));
    CascadeMux I__2136 (
            .O(N__11625),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_ ));
    InMux I__2135 (
            .O(N__11622),
            .I(N__11616));
    InMux I__2134 (
            .O(N__11621),
            .I(N__11616));
    LocalMux I__2133 (
            .O(N__11616),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5 ));
    CascadeMux I__2132 (
            .O(N__11613),
            .I(\Lab_UT.dictrl.un1_state_16_cascade_ ));
    InMux I__2131 (
            .O(N__11610),
            .I(N__11607));
    LocalMux I__2130 (
            .O(N__11607),
            .I(N__11604));
    Span4Mux_h I__2129 (
            .O(N__11604),
            .I(N__11596));
    InMux I__2128 (
            .O(N__11603),
            .I(N__11591));
    InMux I__2127 (
            .O(N__11602),
            .I(N__11591));
    InMux I__2126 (
            .O(N__11601),
            .I(N__11588));
    InMux I__2125 (
            .O(N__11600),
            .I(N__11583));
    InMux I__2124 (
            .O(N__11599),
            .I(N__11583));
    Odrv4 I__2123 (
            .O(N__11596),
            .I(bu_rx_data_5));
    LocalMux I__2122 (
            .O(N__11591),
            .I(bu_rx_data_5));
    LocalMux I__2121 (
            .O(N__11588),
            .I(bu_rx_data_5));
    LocalMux I__2120 (
            .O(N__11583),
            .I(bu_rx_data_5));
    CascadeMux I__2119 (
            .O(N__11574),
            .I(N__11571));
    InMux I__2118 (
            .O(N__11571),
            .I(N__11566));
    InMux I__2117 (
            .O(N__11570),
            .I(N__11563));
    InMux I__2116 (
            .O(N__11569),
            .I(N__11556));
    LocalMux I__2115 (
            .O(N__11566),
            .I(N__11551));
    LocalMux I__2114 (
            .O(N__11563),
            .I(N__11551));
    InMux I__2113 (
            .O(N__11562),
            .I(N__11546));
    InMux I__2112 (
            .O(N__11561),
            .I(N__11546));
    InMux I__2111 (
            .O(N__11560),
            .I(N__11541));
    InMux I__2110 (
            .O(N__11559),
            .I(N__11541));
    LocalMux I__2109 (
            .O(N__11556),
            .I(bu_rx_data_1));
    Odrv4 I__2108 (
            .O(N__11551),
            .I(bu_rx_data_1));
    LocalMux I__2107 (
            .O(N__11546),
            .I(bu_rx_data_1));
    LocalMux I__2106 (
            .O(N__11541),
            .I(bu_rx_data_1));
    InMux I__2105 (
            .O(N__11532),
            .I(N__11525));
    InMux I__2104 (
            .O(N__11531),
            .I(N__11521));
    InMux I__2103 (
            .O(N__11530),
            .I(N__11514));
    InMux I__2102 (
            .O(N__11529),
            .I(N__11514));
    InMux I__2101 (
            .O(N__11528),
            .I(N__11514));
    LocalMux I__2100 (
            .O(N__11525),
            .I(N__11511));
    InMux I__2099 (
            .O(N__11524),
            .I(N__11508));
    LocalMux I__2098 (
            .O(N__11521),
            .I(N__11503));
    LocalMux I__2097 (
            .O(N__11514),
            .I(N__11503));
    Odrv12 I__2096 (
            .O(N__11511),
            .I(bu_rx_data_0));
    LocalMux I__2095 (
            .O(N__11508),
            .I(bu_rx_data_0));
    Odrv4 I__2094 (
            .O(N__11503),
            .I(bu_rx_data_0));
    InMux I__2093 (
            .O(N__11496),
            .I(N__11492));
    InMux I__2092 (
            .O(N__11495),
            .I(N__11489));
    LocalMux I__2091 (
            .O(N__11492),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__2090 (
            .O(N__11489),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__2089 (
            .O(N__11484),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    InMux I__2088 (
            .O(N__11481),
            .I(N__11478));
    LocalMux I__2087 (
            .O(N__11478),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ));
    CascadeMux I__2086 (
            .O(N__11475),
            .I(N__11472));
    InMux I__2085 (
            .O(N__11472),
            .I(N__11469));
    LocalMux I__2084 (
            .O(N__11469),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ));
    InMux I__2083 (
            .O(N__11466),
            .I(N__11462));
    InMux I__2082 (
            .O(N__11465),
            .I(N__11459));
    LocalMux I__2081 (
            .O(N__11462),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__2080 (
            .O(N__11459),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__2079 (
            .O(N__11454),
            .I(N__11451));
    LocalMux I__2078 (
            .O(N__11451),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ));
    CascadeMux I__2077 (
            .O(N__11448),
            .I(N__11444));
    InMux I__2076 (
            .O(N__11447),
            .I(N__11441));
    InMux I__2075 (
            .O(N__11444),
            .I(N__11438));
    LocalMux I__2074 (
            .O(N__11441),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__2073 (
            .O(N__11438),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__2072 (
            .O(N__11433),
            .I(N__11430));
    LocalMux I__2071 (
            .O(N__11430),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_1 ));
    CascadeMux I__2070 (
            .O(N__11427),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_ ));
    CascadeMux I__2069 (
            .O(N__11424),
            .I(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_ ));
    InMux I__2068 (
            .O(N__11421),
            .I(N__11418));
    LocalMux I__2067 (
            .O(N__11418),
            .I(\Lab_UT.dictrl.next_state_out_1 ));
    CascadeMux I__2066 (
            .O(N__11415),
            .I(\Lab_UT.dictrl.N_97_cascade_ ));
    CascadeMux I__2065 (
            .O(N__11412),
            .I(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_ ));
    InMux I__2064 (
            .O(N__11409),
            .I(N__11404));
    InMux I__2063 (
            .O(N__11408),
            .I(N__11401));
    InMux I__2062 (
            .O(N__11407),
            .I(N__11398));
    LocalMux I__2061 (
            .O(N__11404),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__2060 (
            .O(N__11401),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__2059 (
            .O(N__11398),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__2058 (
            .O(N__11391),
            .I(N__11385));
    InMux I__2057 (
            .O(N__11390),
            .I(N__11382));
    InMux I__2056 (
            .O(N__11389),
            .I(N__11379));
    InMux I__2055 (
            .O(N__11388),
            .I(N__11376));
    InMux I__2054 (
            .O(N__11385),
            .I(N__11373));
    LocalMux I__2053 (
            .O(N__11382),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2052 (
            .O(N__11379),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2051 (
            .O(N__11376),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2050 (
            .O(N__11373),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__2049 (
            .O(N__11364),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__2048 (
            .O(N__11361),
            .I(N__11358));
    LocalMux I__2047 (
            .O(N__11358),
            .I(N__11354));
    InMux I__2046 (
            .O(N__11357),
            .I(N__11351));
    Odrv4 I__2045 (
            .O(N__11354),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__2044 (
            .O(N__11351),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__2043 (
            .O(N__11346),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__2042 (
            .O(N__11343),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    CascadeMux I__2041 (
            .O(N__11340),
            .I(\Lab_UT.didp.did_alarmMatch_1_cascade_ ));
    InMux I__2040 (
            .O(N__11337),
            .I(N__11334));
    LocalMux I__2039 (
            .O(N__11334),
            .I(\Lab_UT.zero ));
    InMux I__2038 (
            .O(N__11331),
            .I(N__11325));
    InMux I__2037 (
            .O(N__11330),
            .I(N__11325));
    LocalMux I__2036 (
            .O(N__11325),
            .I(\Lab_UT.alarmMatch ));
    InMux I__2035 (
            .O(N__11322),
            .I(N__11319));
    LocalMux I__2034 (
            .O(N__11319),
            .I(\Lab_UT.didp.countrce3.did_alarmMatch_0 ));
    InMux I__2033 (
            .O(N__11316),
            .I(N__11313));
    LocalMux I__2032 (
            .O(N__11313),
            .I(\Lab_UT.q_5_3 ));
    CascadeMux I__2031 (
            .O(N__11310),
            .I(\Lab_UT.q_5_0_cascade_ ));
    InMux I__2030 (
            .O(N__11307),
            .I(N__11304));
    LocalMux I__2029 (
            .O(N__11304),
            .I(\Lab_UT.q_5_2 ));
    CascadeMux I__2028 (
            .O(N__11301),
            .I(N__11298));
    InMux I__2027 (
            .O(N__11298),
            .I(N__11292));
    InMux I__2026 (
            .O(N__11297),
            .I(N__11292));
    LocalMux I__2025 (
            .O(N__11292),
            .I(N__11289));
    Span4Mux_v I__2024 (
            .O(N__11289),
            .I(N__11286));
    Odrv4 I__2023 (
            .O(N__11286),
            .I(\Lab_UT.N_27_i ));
    InMux I__2022 (
            .O(N__11283),
            .I(N__11280));
    LocalMux I__2021 (
            .O(N__11280),
            .I(N__11277));
    Span4Mux_h I__2020 (
            .O(N__11277),
            .I(N__11274));
    Odrv4 I__2019 (
            .O(N__11274),
            .I(\resetGen.escKeyZ0Z_4 ));
    InMux I__2018 (
            .O(N__11271),
            .I(N__11268));
    LocalMux I__2017 (
            .O(N__11268),
            .I(N__11261));
    InMux I__2016 (
            .O(N__11267),
            .I(N__11252));
    InMux I__2015 (
            .O(N__11266),
            .I(N__11252));
    InMux I__2014 (
            .O(N__11265),
            .I(N__11252));
    InMux I__2013 (
            .O(N__11264),
            .I(N__11252));
    Span4Mux_v I__2012 (
            .O(N__11261),
            .I(N__11247));
    LocalMux I__2011 (
            .O(N__11252),
            .I(N__11247));
    Odrv4 I__2010 (
            .O(N__11247),
            .I(\resetGen.escKeyZ0 ));
    CascadeMux I__2009 (
            .O(N__11244),
            .I(\Lab_UT.bcd2segment1.i2_mux_cascade_ ));
    InMux I__2008 (
            .O(N__11241),
            .I(N__11238));
    LocalMux I__2007 (
            .O(N__11238),
            .I(N__11234));
    InMux I__2006 (
            .O(N__11237),
            .I(N__11231));
    Odrv4 I__2005 (
            .O(N__11234),
            .I(\uu2.bitmapZ0Z_40 ));
    LocalMux I__2004 (
            .O(N__11231),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__2003 (
            .O(N__11226),
            .I(N__11223));
    InMux I__2002 (
            .O(N__11223),
            .I(N__11217));
    InMux I__2001 (
            .O(N__11222),
            .I(N__11217));
    LocalMux I__2000 (
            .O(N__11217),
            .I(\uu2.bitmapZ0Z_296 ));
    CascadeMux I__1999 (
            .O(N__11214),
            .I(\uu2.m95_i_m2_i_m2_1_cascade_ ));
    CascadeMux I__1998 (
            .O(N__11211),
            .I(\uu2.N_16_cascade_ ));
    CascadeMux I__1997 (
            .O(N__11208),
            .I(N__11205));
    InMux I__1996 (
            .O(N__11205),
            .I(N__11200));
    CascadeMux I__1995 (
            .O(N__11204),
            .I(N__11197));
    InMux I__1994 (
            .O(N__11203),
            .I(N__11194));
    LocalMux I__1993 (
            .O(N__11200),
            .I(N__11191));
    InMux I__1992 (
            .O(N__11197),
            .I(N__11188));
    LocalMux I__1991 (
            .O(N__11194),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__1990 (
            .O(N__11191),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__1989 (
            .O(N__11188),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    CascadeMux I__1988 (
            .O(N__11181),
            .I(N__11173));
    CascadeMux I__1987 (
            .O(N__11180),
            .I(N__11169));
    CascadeMux I__1986 (
            .O(N__11179),
            .I(N__11165));
    InMux I__1985 (
            .O(N__11178),
            .I(N__11156));
    InMux I__1984 (
            .O(N__11177),
            .I(N__11156));
    InMux I__1983 (
            .O(N__11176),
            .I(N__11156));
    InMux I__1982 (
            .O(N__11173),
            .I(N__11153));
    InMux I__1981 (
            .O(N__11172),
            .I(N__11142));
    InMux I__1980 (
            .O(N__11169),
            .I(N__11142));
    InMux I__1979 (
            .O(N__11168),
            .I(N__11142));
    InMux I__1978 (
            .O(N__11165),
            .I(N__11142));
    InMux I__1977 (
            .O(N__11164),
            .I(N__11139));
    InMux I__1976 (
            .O(N__11163),
            .I(N__11135));
    LocalMux I__1975 (
            .O(N__11156),
            .I(N__11132));
    LocalMux I__1974 (
            .O(N__11153),
            .I(N__11127));
    InMux I__1973 (
            .O(N__11152),
            .I(N__11122));
    InMux I__1972 (
            .O(N__11151),
            .I(N__11122));
    LocalMux I__1971 (
            .O(N__11142),
            .I(N__11117));
    LocalMux I__1970 (
            .O(N__11139),
            .I(N__11117));
    InMux I__1969 (
            .O(N__11138),
            .I(N__11114));
    LocalMux I__1968 (
            .O(N__11135),
            .I(N__11111));
    Span4Mux_v I__1967 (
            .O(N__11132),
            .I(N__11108));
    InMux I__1966 (
            .O(N__11131),
            .I(N__11103));
    InMux I__1965 (
            .O(N__11130),
            .I(N__11103));
    Span4Mux_h I__1964 (
            .O(N__11127),
            .I(N__11096));
    LocalMux I__1963 (
            .O(N__11122),
            .I(N__11096));
    Span4Mux_h I__1962 (
            .O(N__11117),
            .I(N__11096));
    LocalMux I__1961 (
            .O(N__11114),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1960 (
            .O(N__11111),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1959 (
            .O(N__11108),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1958 (
            .O(N__11103),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1957 (
            .O(N__11096),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    InMux I__1956 (
            .O(N__11085),
            .I(N__11082));
    LocalMux I__1955 (
            .O(N__11082),
            .I(N__11079));
    Odrv4 I__1954 (
            .O(N__11079),
            .I(\uu2.N_67_1_0 ));
    CascadeMux I__1953 (
            .O(N__11076),
            .I(\uu2.N_67_1_0_cascade_ ));
    InMux I__1952 (
            .O(N__11073),
            .I(N__11070));
    LocalMux I__1951 (
            .O(N__11070),
            .I(N__11067));
    Odrv4 I__1950 (
            .O(N__11067),
            .I(\uu2.mem0.N_55_0_0_0 ));
    InMux I__1949 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__1948 (
            .O(N__11061),
            .I(\uu2.mem0.g2_1 ));
    CascadeMux I__1947 (
            .O(N__11058),
            .I(\Lab_UT.bcd2segment1.N_250_cascade_ ));
    InMux I__1946 (
            .O(N__11055),
            .I(N__11052));
    LocalMux I__1945 (
            .O(N__11052),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_34 ));
    InMux I__1944 (
            .O(N__11049),
            .I(N__11046));
    LocalMux I__1943 (
            .O(N__11046),
            .I(N__11043));
    Span4Mux_h I__1942 (
            .O(N__11043),
            .I(N__11038));
    InMux I__1941 (
            .O(N__11042),
            .I(N__11033));
    InMux I__1940 (
            .O(N__11041),
            .I(N__11033));
    Odrv4 I__1939 (
            .O(N__11038),
            .I(L3_tx_data_2));
    LocalMux I__1938 (
            .O(N__11033),
            .I(L3_tx_data_2));
    InMux I__1937 (
            .O(N__11028),
            .I(N__11025));
    LocalMux I__1936 (
            .O(N__11025),
            .I(N__11022));
    Odrv12 I__1935 (
            .O(N__11022),
            .I(\uu2.mem0.N_93_i ));
    InMux I__1934 (
            .O(N__11019),
            .I(N__11016));
    LocalMux I__1933 (
            .O(N__11016),
            .I(\uu2.mem0.N_57_0_0 ));
    InMux I__1932 (
            .O(N__11013),
            .I(N__11010));
    LocalMux I__1931 (
            .O(N__11010),
            .I(\uu2.mem0.N_67_0 ));
    CascadeMux I__1930 (
            .O(N__11007),
            .I(\uu2.mem0.g0_1_cascade_ ));
    InMux I__1929 (
            .O(N__11004),
            .I(N__11001));
    LocalMux I__1928 (
            .O(N__11001),
            .I(\uu2.mem0.g0_2 ));
    InMux I__1927 (
            .O(N__10998),
            .I(N__10995));
    LocalMux I__1926 (
            .O(N__10995),
            .I(\uu2.mem0.i14_mux ));
    InMux I__1925 (
            .O(N__10992),
            .I(N__10989));
    LocalMux I__1924 (
            .O(N__10989),
            .I(N__10986));
    Span4Mux_h I__1923 (
            .O(N__10986),
            .I(N__10983));
    Odrv4 I__1922 (
            .O(N__10983),
            .I(\uu2.mem0.N_126_0 ));
    CascadeMux I__1921 (
            .O(N__10980),
            .I(\uu2.mem0.g0_1_3_cascade_ ));
    InMux I__1920 (
            .O(N__10977),
            .I(N__10974));
    LocalMux I__1919 (
            .O(N__10974),
            .I(\uu2.mem0.G_13_0_a2_0_1 ));
    CascadeMux I__1918 (
            .O(N__10971),
            .I(\uu2.mem0.N_22_cascade_ ));
    InMux I__1917 (
            .O(N__10968),
            .I(N__10965));
    LocalMux I__1916 (
            .O(N__10965),
            .I(N__10962));
    Span4Mux_h I__1915 (
            .O(N__10962),
            .I(N__10959));
    Odrv4 I__1914 (
            .O(N__10959),
            .I(\uu2.mem0.N_66_0_i ));
    InMux I__1913 (
            .O(N__10956),
            .I(N__10953));
    LocalMux I__1912 (
            .O(N__10953),
            .I(\uu2.mem0.g0_i_m2_1 ));
    InMux I__1911 (
            .O(N__10950),
            .I(N__10947));
    LocalMux I__1910 (
            .O(N__10947),
            .I(N__10944));
    Span4Mux_h I__1909 (
            .O(N__10944),
            .I(N__10941));
    Odrv4 I__1908 (
            .O(N__10941),
            .I(\uu2.mem0.g2_0_0_0 ));
    CascadeMux I__1907 (
            .O(N__10938),
            .I(N__10935));
    InMux I__1906 (
            .O(N__10935),
            .I(N__10932));
    LocalMux I__1905 (
            .O(N__10932),
            .I(\uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1 ));
    CascadeMux I__1904 (
            .O(N__10929),
            .I(\uu2.mem0.N_92_0_cascade_ ));
    InMux I__1903 (
            .O(N__10926),
            .I(N__10923));
    LocalMux I__1902 (
            .O(N__10923),
            .I(\uu2.mem0.m73_ns_1_0 ));
    InMux I__1901 (
            .O(N__10920),
            .I(N__10917));
    LocalMux I__1900 (
            .O(N__10917),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_1_4 ));
    CascadeMux I__1899 (
            .O(N__10914),
            .I(N__10911));
    InMux I__1898 (
            .O(N__10911),
            .I(N__10905));
    InMux I__1897 (
            .O(N__10910),
            .I(N__10905));
    LocalMux I__1896 (
            .O(N__10905),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__1895 (
            .O(N__10902),
            .I(N__10896));
    InMux I__1894 (
            .O(N__10901),
            .I(N__10896));
    LocalMux I__1893 (
            .O(N__10896),
            .I(\uu2.bitmapZ0Z_90 ));
    CascadeMux I__1892 (
            .O(N__10893),
            .I(\uu2.mem0.N_92_0_0_cascade_ ));
    CascadeMux I__1891 (
            .O(N__10890),
            .I(N__10887));
    InMux I__1890 (
            .O(N__10887),
            .I(N__10884));
    LocalMux I__1889 (
            .O(N__10884),
            .I(N__10881));
    Odrv4 I__1888 (
            .O(N__10881),
            .I(\uu2.mem0.m73_ns_1_0_0_1 ));
    InMux I__1887 (
            .O(N__10878),
            .I(N__10875));
    LocalMux I__1886 (
            .O(N__10875),
            .I(\uu2.mem0.N_74_0 ));
    InMux I__1885 (
            .O(N__10872),
            .I(N__10869));
    LocalMux I__1884 (
            .O(N__10869),
            .I(N__10866));
    Odrv4 I__1883 (
            .O(N__10866),
            .I(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0 ));
    CascadeMux I__1882 (
            .O(N__10863),
            .I(\Lab_UT.bcd2segment1.N_194_cascade_ ));
    CascadeMux I__1881 (
            .O(N__10860),
            .I(\buart.Z_rx.ser_clk_2_cascade_ ));
    CascadeMux I__1880 (
            .O(N__10857),
            .I(\Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_ ));
    CascadeMux I__1879 (
            .O(N__10854),
            .I(N__10851));
    InMux I__1878 (
            .O(N__10851),
            .I(N__10848));
    LocalMux I__1877 (
            .O(N__10848),
            .I(N__10843));
    InMux I__1876 (
            .O(N__10847),
            .I(N__10840));
    InMux I__1875 (
            .O(N__10846),
            .I(N__10837));
    Span4Mux_h I__1874 (
            .O(N__10843),
            .I(N__10834));
    LocalMux I__1873 (
            .O(N__10840),
            .I(N__10829));
    LocalMux I__1872 (
            .O(N__10837),
            .I(N__10829));
    Odrv4 I__1871 (
            .O(N__10834),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z4 ));
    Odrv4 I__1870 (
            .O(N__10829),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z4 ));
    InMux I__1869 (
            .O(N__10824),
            .I(N__10821));
    LocalMux I__1868 (
            .O(N__10821),
            .I(\Lab_UT.dictrl.next_alarmstate4Z0Z_0 ));
    CascadeMux I__1867 (
            .O(N__10818),
            .I(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_ ));
    CascadeMux I__1866 (
            .O(N__10815),
            .I(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ));
    CascadeMux I__1865 (
            .O(N__10812),
            .I(\Lab_UT.bcd2segment1.N_222_cascade_ ));
    InMux I__1864 (
            .O(N__10809),
            .I(N__10804));
    InMux I__1863 (
            .O(N__10808),
            .I(N__10798));
    InMux I__1862 (
            .O(N__10807),
            .I(N__10795));
    LocalMux I__1861 (
            .O(N__10804),
            .I(N__10792));
    InMux I__1860 (
            .O(N__10803),
            .I(N__10785));
    InMux I__1859 (
            .O(N__10802),
            .I(N__10785));
    InMux I__1858 (
            .O(N__10801),
            .I(N__10785));
    LocalMux I__1857 (
            .O(N__10798),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    LocalMux I__1856 (
            .O(N__10795),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    Odrv4 I__1855 (
            .O(N__10792),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    LocalMux I__1854 (
            .O(N__10785),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    InMux I__1853 (
            .O(N__10776),
            .I(N__10773));
    LocalMux I__1852 (
            .O(N__10773),
            .I(N__10767));
    InMux I__1851 (
            .O(N__10772),
            .I(N__10764));
    InMux I__1850 (
            .O(N__10771),
            .I(N__10759));
    InMux I__1849 (
            .O(N__10770),
            .I(N__10759));
    Odrv4 I__1848 (
            .O(N__10767),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__1847 (
            .O(N__10764),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__1846 (
            .O(N__10759),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    InMux I__1845 (
            .O(N__10752),
            .I(N__10748));
    InMux I__1844 (
            .O(N__10751),
            .I(N__10745));
    LocalMux I__1843 (
            .O(N__10748),
            .I(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ));
    LocalMux I__1842 (
            .O(N__10745),
            .I(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ));
    InMux I__1841 (
            .O(N__10740),
            .I(N__10735));
    InMux I__1840 (
            .O(N__10739),
            .I(N__10732));
    InMux I__1839 (
            .O(N__10738),
            .I(N__10729));
    LocalMux I__1838 (
            .O(N__10735),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__1837 (
            .O(N__10732),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__1836 (
            .O(N__10729),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__1835 (
            .O(N__10722),
            .I(N__10718));
    InMux I__1834 (
            .O(N__10721),
            .I(N__10712));
    LocalMux I__1833 (
            .O(N__10718),
            .I(N__10709));
    InMux I__1832 (
            .O(N__10717),
            .I(N__10702));
    InMux I__1831 (
            .O(N__10716),
            .I(N__10702));
    InMux I__1830 (
            .O(N__10715),
            .I(N__10702));
    LocalMux I__1829 (
            .O(N__10712),
            .I(\uu2.l_countZ0Z_4 ));
    Odrv4 I__1828 (
            .O(N__10709),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__1827 (
            .O(N__10702),
            .I(\uu2.l_countZ0Z_4 ));
    CascadeMux I__1826 (
            .O(N__10695),
            .I(N__10691));
    InMux I__1825 (
            .O(N__10694),
            .I(N__10686));
    InMux I__1824 (
            .O(N__10691),
            .I(N__10686));
    LocalMux I__1823 (
            .O(N__10686),
            .I(N__10682));
    InMux I__1822 (
            .O(N__10685),
            .I(N__10679));
    Span4Mux_v I__1821 (
            .O(N__10682),
            .I(N__10676));
    LocalMux I__1820 (
            .O(N__10679),
            .I(N__10671));
    Sp12to4 I__1819 (
            .O(N__10676),
            .I(N__10671));
    Odrv12 I__1818 (
            .O(N__10671),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    CascadeMux I__1817 (
            .O(N__10668),
            .I(\Lab_UT.q_5_1_cascade_ ));
    CascadeMux I__1816 (
            .O(N__10665),
            .I(\Lab_UT.bcd2segment1.i5_mux_cascade_ ));
    InMux I__1815 (
            .O(N__10662),
            .I(N__10653));
    InMux I__1814 (
            .O(N__10661),
            .I(N__10648));
    InMux I__1813 (
            .O(N__10660),
            .I(N__10648));
    InMux I__1812 (
            .O(N__10659),
            .I(N__10645));
    InMux I__1811 (
            .O(N__10658),
            .I(N__10640));
    InMux I__1810 (
            .O(N__10657),
            .I(N__10640));
    CascadeMux I__1809 (
            .O(N__10656),
            .I(N__10636));
    LocalMux I__1808 (
            .O(N__10653),
            .I(N__10631));
    LocalMux I__1807 (
            .O(N__10648),
            .I(N__10624));
    LocalMux I__1806 (
            .O(N__10645),
            .I(N__10624));
    LocalMux I__1805 (
            .O(N__10640),
            .I(N__10624));
    InMux I__1804 (
            .O(N__10639),
            .I(N__10617));
    InMux I__1803 (
            .O(N__10636),
            .I(N__10617));
    InMux I__1802 (
            .O(N__10635),
            .I(N__10617));
    InMux I__1801 (
            .O(N__10634),
            .I(N__10614));
    Span4Mux_v I__1800 (
            .O(N__10631),
            .I(N__10611));
    Span4Mux_v I__1799 (
            .O(N__10624),
            .I(N__10608));
    LocalMux I__1798 (
            .O(N__10617),
            .I(\Lab_UT.cnt_2 ));
    LocalMux I__1797 (
            .O(N__10614),
            .I(\Lab_UT.cnt_2 ));
    Odrv4 I__1796 (
            .O(N__10611),
            .I(\Lab_UT.cnt_2 ));
    Odrv4 I__1795 (
            .O(N__10608),
            .I(\Lab_UT.cnt_2 ));
    CascadeMux I__1794 (
            .O(N__10599),
            .I(\Lab_UT.bcd2segment1.m42_amZ0_cascade_ ));
    InMux I__1793 (
            .O(N__10596),
            .I(N__10593));
    LocalMux I__1792 (
            .O(N__10593),
            .I(\Lab_UT.bcd2segment1.m52_bmZ0 ));
    InMux I__1791 (
            .O(N__10590),
            .I(N__10587));
    LocalMux I__1790 (
            .O(N__10587),
            .I(\Lab_UT.bcd2segment1.N_42_i ));
    InMux I__1789 (
            .O(N__10584),
            .I(N__10579));
    InMux I__1788 (
            .O(N__10583),
            .I(N__10576));
    InMux I__1787 (
            .O(N__10582),
            .I(N__10573));
    LocalMux I__1786 (
            .O(N__10579),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_0 ));
    LocalMux I__1785 (
            .O(N__10576),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_0 ));
    LocalMux I__1784 (
            .O(N__10573),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_0 ));
    CascadeMux I__1783 (
            .O(N__10566),
            .I(\Lab_UT.dictrl.idle_cascade_ ));
    InMux I__1782 (
            .O(N__10563),
            .I(N__10556));
    InMux I__1781 (
            .O(N__10562),
            .I(N__10556));
    InMux I__1780 (
            .O(N__10561),
            .I(N__10553));
    LocalMux I__1779 (
            .O(N__10556),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    LocalMux I__1778 (
            .O(N__10553),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    CascadeMux I__1777 (
            .O(N__10548),
            .I(N__10545));
    InMux I__1776 (
            .O(N__10545),
            .I(N__10542));
    LocalMux I__1775 (
            .O(N__10542),
            .I(N__10539));
    Span4Mux_h I__1774 (
            .O(N__10539),
            .I(N__10536));
    Odrv4 I__1773 (
            .O(N__10536),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_0 ));
    IoInMux I__1772 (
            .O(N__10533),
            .I(N__10529));
    InMux I__1771 (
            .O(N__10532),
            .I(N__10526));
    LocalMux I__1770 (
            .O(N__10529),
            .I(N__10523));
    LocalMux I__1769 (
            .O(N__10526),
            .I(N__10520));
    Span12Mux_s9_v I__1768 (
            .O(N__10523),
            .I(N__10517));
    Span4Mux_v I__1767 (
            .O(N__10520),
            .I(N__10514));
    Odrv12 I__1766 (
            .O(N__10517),
            .I(clk));
    Odrv4 I__1765 (
            .O(N__10514),
            .I(clk));
    SRMux I__1764 (
            .O(N__10509),
            .I(N__10505));
    CEMux I__1763 (
            .O(N__10508),
            .I(N__10502));
    LocalMux I__1762 (
            .O(N__10505),
            .I(N__10499));
    LocalMux I__1761 (
            .O(N__10502),
            .I(N__10496));
    Span4Mux_h I__1760 (
            .O(N__10499),
            .I(N__10491));
    Span4Mux_h I__1759 (
            .O(N__10496),
            .I(N__10491));
    Odrv4 I__1758 (
            .O(N__10491),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1757 (
            .O(N__10488),
            .I(\uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_ ));
    InMux I__1756 (
            .O(N__10485),
            .I(N__10482));
    LocalMux I__1755 (
            .O(N__10482),
            .I(N__10479));
    Span4Mux_h I__1754 (
            .O(N__10479),
            .I(N__10476));
    Odrv4 I__1753 (
            .O(N__10476),
            .I(\uu2.mem0.g1_2_0 ));
    InMux I__1752 (
            .O(N__10473),
            .I(N__10470));
    LocalMux I__1751 (
            .O(N__10470),
            .I(\uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0 ));
    InMux I__1750 (
            .O(N__10467),
            .I(N__10464));
    LocalMux I__1749 (
            .O(N__10464),
            .I(\uu2.mem0.g0_7_0_0_1 ));
    CascadeMux I__1748 (
            .O(N__10461),
            .I(\Lab_UT.alarmchar9_cascade_ ));
    InMux I__1747 (
            .O(N__10458),
            .I(N__10455));
    LocalMux I__1746 (
            .O(N__10455),
            .I(N__10452));
    Span4Mux_h I__1745 (
            .O(N__10452),
            .I(N__10449));
    Odrv4 I__1744 (
            .O(N__10449),
            .I(\Lab_UT.alarmcharZ0Z_2 ));
    InMux I__1743 (
            .O(N__10446),
            .I(N__10443));
    LocalMux I__1742 (
            .O(N__10443),
            .I(\Lab_UT.bcd2segment1.N_160 ));
    CascadeMux I__1741 (
            .O(N__10440),
            .I(\uu2.mem0.N_3_0_cascade_ ));
    InMux I__1740 (
            .O(N__10437),
            .I(N__10434));
    LocalMux I__1739 (
            .O(N__10434),
            .I(\uu2.mem0.N_98_0_0_0 ));
    InMux I__1738 (
            .O(N__10431),
            .I(N__10426));
    InMux I__1737 (
            .O(N__10430),
            .I(N__10423));
    InMux I__1736 (
            .O(N__10429),
            .I(N__10420));
    LocalMux I__1735 (
            .O(N__10426),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    LocalMux I__1734 (
            .O(N__10423),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    LocalMux I__1733 (
            .O(N__10420),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    InMux I__1732 (
            .O(N__10413),
            .I(N__10407));
    InMux I__1731 (
            .O(N__10412),
            .I(N__10407));
    LocalMux I__1730 (
            .O(N__10407),
            .I(\uu2.N_1585_0_0 ));
    CascadeMux I__1729 (
            .O(N__10404),
            .I(\Lab_UT.bcd2segment1.i6_mux_cascade_ ));
    InMux I__1728 (
            .O(N__10401),
            .I(N__10398));
    LocalMux I__1727 (
            .O(N__10398),
            .I(\Lab_UT.bcd2segment1.m68_amZ0 ));
    InMux I__1726 (
            .O(N__10395),
            .I(N__10392));
    LocalMux I__1725 (
            .O(N__10392),
            .I(N__10384));
    InMux I__1724 (
            .O(N__10391),
            .I(N__10375));
    InMux I__1723 (
            .O(N__10390),
            .I(N__10375));
    InMux I__1722 (
            .O(N__10389),
            .I(N__10375));
    InMux I__1721 (
            .O(N__10388),
            .I(N__10375));
    InMux I__1720 (
            .O(N__10387),
            .I(N__10372));
    Span4Mux_h I__1719 (
            .O(N__10384),
            .I(N__10369));
    LocalMux I__1718 (
            .O(N__10375),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__1717 (
            .O(N__10372),
            .I(\resetGen.reset_countZ0Z_4 ));
    Odrv4 I__1716 (
            .O(N__10369),
            .I(\resetGen.reset_countZ0Z_4 ));
    IoInMux I__1715 (
            .O(N__10362),
            .I(N__10359));
    LocalMux I__1714 (
            .O(N__10359),
            .I(N__10354));
    InMux I__1713 (
            .O(N__10358),
            .I(N__10351));
    InMux I__1712 (
            .O(N__10357),
            .I(N__10346));
    IoSpan4Mux I__1711 (
            .O(N__10354),
            .I(N__10343));
    LocalMux I__1710 (
            .O(N__10351),
            .I(N__10340));
    InMux I__1709 (
            .O(N__10350),
            .I(N__10334));
    InMux I__1708 (
            .O(N__10349),
            .I(N__10334));
    LocalMux I__1707 (
            .O(N__10346),
            .I(N__10329));
    Span4Mux_s1_h I__1706 (
            .O(N__10343),
            .I(N__10329));
    Span4Mux_v I__1705 (
            .O(N__10340),
            .I(N__10326));
    InMux I__1704 (
            .O(N__10339),
            .I(N__10323));
    LocalMux I__1703 (
            .O(N__10334),
            .I(N__10318));
    Span4Mux_h I__1702 (
            .O(N__10329),
            .I(N__10318));
    Odrv4 I__1701 (
            .O(N__10326),
            .I(rst));
    LocalMux I__1700 (
            .O(N__10323),
            .I(rst));
    Odrv4 I__1699 (
            .O(N__10318),
            .I(rst));
    CascadeMux I__1698 (
            .O(N__10311),
            .I(N__10307));
    InMux I__1697 (
            .O(N__10310),
            .I(N__10302));
    InMux I__1696 (
            .O(N__10307),
            .I(N__10298));
    InMux I__1695 (
            .O(N__10306),
            .I(N__10295));
    CascadeMux I__1694 (
            .O(N__10305),
            .I(N__10292));
    LocalMux I__1693 (
            .O(N__10302),
            .I(N__10289));
    InMux I__1692 (
            .O(N__10301),
            .I(N__10286));
    LocalMux I__1691 (
            .O(N__10298),
            .I(N__10283));
    LocalMux I__1690 (
            .O(N__10295),
            .I(N__10280));
    InMux I__1689 (
            .O(N__10292),
            .I(N__10277));
    Span4Mux_v I__1688 (
            .O(N__10289),
            .I(N__10274));
    LocalMux I__1687 (
            .O(N__10286),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1686 (
            .O(N__10283),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1685 (
            .O(N__10280),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__1684 (
            .O(N__10277),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1683 (
            .O(N__10274),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__1682 (
            .O(N__10263),
            .I(\uu2.mem0.N_17_0_cascade_ ));
    CascadeMux I__1681 (
            .O(N__10260),
            .I(N__10257));
    InMux I__1680 (
            .O(N__10257),
            .I(N__10252));
    CascadeMux I__1679 (
            .O(N__10256),
            .I(N__10246));
    CascadeMux I__1678 (
            .O(N__10255),
            .I(N__10243));
    LocalMux I__1677 (
            .O(N__10252),
            .I(N__10240));
    CascadeMux I__1676 (
            .O(N__10251),
            .I(N__10237));
    InMux I__1675 (
            .O(N__10250),
            .I(N__10230));
    InMux I__1674 (
            .O(N__10249),
            .I(N__10230));
    InMux I__1673 (
            .O(N__10246),
            .I(N__10230));
    InMux I__1672 (
            .O(N__10243),
            .I(N__10227));
    Span4Mux_v I__1671 (
            .O(N__10240),
            .I(N__10224));
    InMux I__1670 (
            .O(N__10237),
            .I(N__10221));
    LocalMux I__1669 (
            .O(N__10230),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__1668 (
            .O(N__10227),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__1667 (
            .O(N__10224),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__1666 (
            .O(N__10221),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__1665 (
            .O(N__10212),
            .I(N__10209));
    InMux I__1664 (
            .O(N__10209),
            .I(N__10206));
    LocalMux I__1663 (
            .O(N__10206),
            .I(N__10203));
    Odrv4 I__1662 (
            .O(N__10203),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_5 ));
    InMux I__1661 (
            .O(N__10200),
            .I(N__10197));
    LocalMux I__1660 (
            .O(N__10197),
            .I(N__10194));
    Odrv4 I__1659 (
            .O(N__10194),
            .I(\uu2.mem0.N_107_0_0 ));
    CascadeMux I__1658 (
            .O(N__10191),
            .I(N__10188));
    InMux I__1657 (
            .O(N__10188),
            .I(N__10185));
    LocalMux I__1656 (
            .O(N__10185),
            .I(\uu2.mem0.N_74_0_0_1 ));
    CascadeMux I__1655 (
            .O(N__10182),
            .I(\uu2.mem0.g0_7_0_0_2_cascade_ ));
    CascadeMux I__1654 (
            .O(N__10179),
            .I(\Lab_UT.bcd2segment1.N_187_cascade_ ));
    CascadeMux I__1653 (
            .O(N__10176),
            .I(\Lab_UT.bcd2segment1.N_189_cascade_ ));
    InMux I__1652 (
            .O(N__10173),
            .I(N__10167));
    InMux I__1651 (
            .O(N__10172),
            .I(N__10167));
    LocalMux I__1650 (
            .O(N__10167),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__1649 (
            .O(N__10164),
            .I(N__10161));
    InMux I__1648 (
            .O(N__10161),
            .I(N__10155));
    InMux I__1647 (
            .O(N__10160),
            .I(N__10155));
    LocalMux I__1646 (
            .O(N__10155),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__1645 (
            .O(N__10152),
            .I(\uu2.mem0.N_107_0_cascade_ ));
    InMux I__1644 (
            .O(N__10149),
            .I(N__10143));
    InMux I__1643 (
            .O(N__10148),
            .I(N__10140));
    InMux I__1642 (
            .O(N__10147),
            .I(N__10135));
    InMux I__1641 (
            .O(N__10146),
            .I(N__10135));
    LocalMux I__1640 (
            .O(N__10143),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1639 (
            .O(N__10140),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1638 (
            .O(N__10135),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__1637 (
            .O(N__10128),
            .I(N__10125));
    InMux I__1636 (
            .O(N__10125),
            .I(N__10122));
    LocalMux I__1635 (
            .O(N__10122),
            .I(N__10119));
    Span4Mux_s3_h I__1634 (
            .O(N__10119),
            .I(N__10116));
    Odrv4 I__1633 (
            .O(N__10116),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_1 ));
    InMux I__1632 (
            .O(N__10113),
            .I(N__10110));
    LocalMux I__1631 (
            .O(N__10110),
            .I(N__10106));
    CascadeMux I__1630 (
            .O(N__10109),
            .I(N__10102));
    Span4Mux_v I__1629 (
            .O(N__10106),
            .I(N__10099));
    InMux I__1628 (
            .O(N__10105),
            .I(N__10094));
    InMux I__1627 (
            .O(N__10102),
            .I(N__10094));
    Odrv4 I__1626 (
            .O(N__10099),
            .I(L3_tx_data_6));
    LocalMux I__1625 (
            .O(N__10094),
            .I(L3_tx_data_6));
    CascadeMux I__1624 (
            .O(N__10089),
            .I(\uu2.mem0.N_130_mux_cascade_ ));
    InMux I__1623 (
            .O(N__10086),
            .I(N__10083));
    LocalMux I__1622 (
            .O(N__10083),
            .I(N__10080));
    Span4Mux_h I__1621 (
            .O(N__10080),
            .I(N__10077));
    Odrv4 I__1620 (
            .O(N__10077),
            .I(\uu2.mem0.N_54_0_i ));
    InMux I__1619 (
            .O(N__10074),
            .I(N__10070));
    InMux I__1618 (
            .O(N__10073),
            .I(N__10066));
    LocalMux I__1617 (
            .O(N__10070),
            .I(N__10063));
    InMux I__1616 (
            .O(N__10069),
            .I(N__10060));
    LocalMux I__1615 (
            .O(N__10066),
            .I(N__10052));
    Span4Mux_v I__1614 (
            .O(N__10063),
            .I(N__10052));
    LocalMux I__1613 (
            .O(N__10060),
            .I(N__10052));
    InMux I__1612 (
            .O(N__10059),
            .I(N__10049));
    Span4Mux_h I__1611 (
            .O(N__10052),
            .I(N__10046));
    LocalMux I__1610 (
            .O(N__10049),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__1609 (
            .O(N__10046),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__1608 (
            .O(N__10041),
            .I(N__10036));
    InMux I__1607 (
            .O(N__10040),
            .I(N__10031));
    InMux I__1606 (
            .O(N__10039),
            .I(N__10031));
    LocalMux I__1605 (
            .O(N__10036),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__1604 (
            .O(N__10031),
            .I(\uu2.un1_l_count_2_0 ));
    InMux I__1603 (
            .O(N__10026),
            .I(N__10021));
    InMux I__1602 (
            .O(N__10025),
            .I(N__10016));
    InMux I__1601 (
            .O(N__10024),
            .I(N__10016));
    LocalMux I__1600 (
            .O(N__10021),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__1599 (
            .O(N__10016),
            .I(\uu2.l_countZ0Z_3 ));
    InMux I__1598 (
            .O(N__10011),
            .I(N__10008));
    LocalMux I__1597 (
            .O(N__10008),
            .I(N__10004));
    InMux I__1596 (
            .O(N__10007),
            .I(N__10001));
    Odrv4 I__1595 (
            .O(N__10004),
            .I(\uu0.delay_lineZ0Z_0 ));
    LocalMux I__1594 (
            .O(N__10001),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__1593 (
            .O(N__9996),
            .I(N__9993));
    LocalMux I__1592 (
            .O(N__9993),
            .I(N__9990));
    Span4Mux_h I__1591 (
            .O(N__9990),
            .I(N__9987));
    Odrv4 I__1590 (
            .O(N__9987),
            .I(\uu0.delay_lineZ0Z_1 ));
    CascadeMux I__1589 (
            .O(N__9984),
            .I(N__9981));
    InMux I__1588 (
            .O(N__9981),
            .I(N__9977));
    InMux I__1587 (
            .O(N__9980),
            .I(N__9974));
    LocalMux I__1586 (
            .O(N__9977),
            .I(\uu2.un284_ci ));
    LocalMux I__1585 (
            .O(N__9974),
            .I(\uu2.un284_ci ));
    CascadeMux I__1584 (
            .O(N__9969),
            .I(N__9962));
    InMux I__1583 (
            .O(N__9968),
            .I(N__9959));
    InMux I__1582 (
            .O(N__9967),
            .I(N__9956));
    InMux I__1581 (
            .O(N__9966),
            .I(N__9951));
    InMux I__1580 (
            .O(N__9965),
            .I(N__9951));
    InMux I__1579 (
            .O(N__9962),
            .I(N__9948));
    LocalMux I__1578 (
            .O(N__9959),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__1577 (
            .O(N__9956),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__1576 (
            .O(N__9951),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__1575 (
            .O(N__9948),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__1574 (
            .O(N__9939),
            .I(N__9936));
    LocalMux I__1573 (
            .O(N__9936),
            .I(N__9933));
    Span4Mux_h I__1572 (
            .O(N__9933),
            .I(N__9930));
    IoSpan4Mux I__1571 (
            .O(N__9930),
            .I(N__9927));
    Odrv4 I__1570 (
            .O(N__9927),
            .I(uart_RXD));
    InMux I__1569 (
            .O(N__9924),
            .I(N__9920));
    InMux I__1568 (
            .O(N__9923),
            .I(N__9917));
    LocalMux I__1567 (
            .O(N__9920),
            .I(N__9914));
    LocalMux I__1566 (
            .O(N__9917),
            .I(\uu2.un350_ci ));
    Odrv4 I__1565 (
            .O(N__9914),
            .I(\uu2.un350_ci ));
    CascadeMux I__1564 (
            .O(N__9909),
            .I(N__9904));
    InMux I__1563 (
            .O(N__9908),
            .I(N__9901));
    InMux I__1562 (
            .O(N__9907),
            .I(N__9898));
    InMux I__1561 (
            .O(N__9904),
            .I(N__9895));
    LocalMux I__1560 (
            .O(N__9901),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1559 (
            .O(N__9898),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1558 (
            .O(N__9895),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__1557 (
            .O(N__9888),
            .I(N__9885));
    InMux I__1556 (
            .O(N__9885),
            .I(N__9880));
    InMux I__1555 (
            .O(N__9884),
            .I(N__9875));
    InMux I__1554 (
            .O(N__9883),
            .I(N__9875));
    LocalMux I__1553 (
            .O(N__9880),
            .I(N__9868));
    LocalMux I__1552 (
            .O(N__9875),
            .I(N__9868));
    InMux I__1551 (
            .O(N__9874),
            .I(N__9863));
    InMux I__1550 (
            .O(N__9873),
            .I(N__9863));
    Span4Mux_h I__1549 (
            .O(N__9868),
            .I(N__9860));
    LocalMux I__1548 (
            .O(N__9863),
            .I(N__9857));
    Odrv4 I__1547 (
            .O(N__9860),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    Odrv12 I__1546 (
            .O(N__9857),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    CEMux I__1545 (
            .O(N__9852),
            .I(N__9849));
    LocalMux I__1544 (
            .O(N__9849),
            .I(N__9846));
    Sp12to4 I__1543 (
            .O(N__9846),
            .I(N__9843));
    Odrv12 I__1542 (
            .O(N__9843),
            .I(\Lab_UT.dictrl.G_74 ));
    InMux I__1541 (
            .O(N__9840),
            .I(N__9833));
    InMux I__1540 (
            .O(N__9839),
            .I(N__9833));
    InMux I__1539 (
            .O(N__9838),
            .I(N__9830));
    LocalMux I__1538 (
            .O(N__9833),
            .I(N__9822));
    LocalMux I__1537 (
            .O(N__9830),
            .I(N__9822));
    InMux I__1536 (
            .O(N__9829),
            .I(N__9815));
    InMux I__1535 (
            .O(N__9828),
            .I(N__9815));
    InMux I__1534 (
            .O(N__9827),
            .I(N__9815));
    Odrv4 I__1533 (
            .O(N__9822),
            .I(\Lab_UT.dictrl.un1_next_alarmstate21_0 ));
    LocalMux I__1532 (
            .O(N__9815),
            .I(\Lab_UT.dictrl.un1_next_alarmstate21_0 ));
    InMux I__1531 (
            .O(N__9810),
            .I(N__9806));
    InMux I__1530 (
            .O(N__9809),
            .I(N__9803));
    LocalMux I__1529 (
            .O(N__9806),
            .I(N__9798));
    LocalMux I__1528 (
            .O(N__9803),
            .I(N__9798));
    Span12Mux_s9_v I__1527 (
            .O(N__9798),
            .I(N__9792));
    InMux I__1526 (
            .O(N__9797),
            .I(N__9785));
    InMux I__1525 (
            .O(N__9796),
            .I(N__9785));
    InMux I__1524 (
            .O(N__9795),
            .I(N__9785));
    Odrv12 I__1523 (
            .O(N__9792),
            .I(\Lab_UT.cnt_0 ));
    LocalMux I__1522 (
            .O(N__9785),
            .I(\Lab_UT.cnt_0 ));
    InMux I__1521 (
            .O(N__9780),
            .I(N__9771));
    InMux I__1520 (
            .O(N__9779),
            .I(N__9771));
    InMux I__1519 (
            .O(N__9778),
            .I(N__9768));
    InMux I__1518 (
            .O(N__9777),
            .I(N__9763));
    InMux I__1517 (
            .O(N__9776),
            .I(N__9763));
    LocalMux I__1516 (
            .O(N__9771),
            .I(N__9760));
    LocalMux I__1515 (
            .O(N__9768),
            .I(\uu2.un306_ci ));
    LocalMux I__1514 (
            .O(N__9763),
            .I(\uu2.un306_ci ));
    Odrv4 I__1513 (
            .O(N__9760),
            .I(\uu2.un306_ci ));
    InMux I__1512 (
            .O(N__9753),
            .I(N__9750));
    LocalMux I__1511 (
            .O(N__9750),
            .I(N__9743));
    InMux I__1510 (
            .O(N__9749),
            .I(N__9738));
    InMux I__1509 (
            .O(N__9748),
            .I(N__9738));
    InMux I__1508 (
            .O(N__9747),
            .I(N__9733));
    InMux I__1507 (
            .O(N__9746),
            .I(N__9733));
    Odrv4 I__1506 (
            .O(N__9743),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__1505 (
            .O(N__9738),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__1504 (
            .O(N__9733),
            .I(\uu2.l_countZ0Z_6 ));
    InMux I__1503 (
            .O(N__9726),
            .I(N__9723));
    LocalMux I__1502 (
            .O(N__9723),
            .I(N__9716));
    InMux I__1501 (
            .O(N__9722),
            .I(N__9709));
    InMux I__1500 (
            .O(N__9721),
            .I(N__9709));
    InMux I__1499 (
            .O(N__9720),
            .I(N__9709));
    InMux I__1498 (
            .O(N__9719),
            .I(N__9706));
    Span4Mux_h I__1497 (
            .O(N__9716),
            .I(N__9696));
    LocalMux I__1496 (
            .O(N__9709),
            .I(N__9691));
    LocalMux I__1495 (
            .O(N__9706),
            .I(N__9691));
    InMux I__1494 (
            .O(N__9705),
            .I(N__9686));
    InMux I__1493 (
            .O(N__9704),
            .I(N__9686));
    InMux I__1492 (
            .O(N__9703),
            .I(N__9679));
    InMux I__1491 (
            .O(N__9702),
            .I(N__9679));
    InMux I__1490 (
            .O(N__9701),
            .I(N__9679));
    InMux I__1489 (
            .O(N__9700),
            .I(N__9674));
    InMux I__1488 (
            .O(N__9699),
            .I(N__9674));
    Odrv4 I__1487 (
            .O(N__9696),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1486 (
            .O(N__9691),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1485 (
            .O(N__9686),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1484 (
            .O(N__9679),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1483 (
            .O(N__9674),
            .I(\uu0.un4_l_count_0 ));
    InMux I__1482 (
            .O(N__9663),
            .I(N__9660));
    LocalMux I__1481 (
            .O(N__9660),
            .I(N__9656));
    InMux I__1480 (
            .O(N__9659),
            .I(N__9653));
    Span4Mux_v I__1479 (
            .O(N__9656),
            .I(N__9647));
    LocalMux I__1478 (
            .O(N__9653),
            .I(N__9647));
    InMux I__1477 (
            .O(N__9652),
            .I(N__9644));
    Span4Mux_v I__1476 (
            .O(N__9647),
            .I(N__9638));
    LocalMux I__1475 (
            .O(N__9644),
            .I(N__9638));
    InMux I__1474 (
            .O(N__9643),
            .I(N__9635));
    Span4Mux_v I__1473 (
            .O(N__9638),
            .I(N__9632));
    LocalMux I__1472 (
            .O(N__9635),
            .I(o_One_Sec_Pulse));
    Odrv4 I__1471 (
            .O(N__9632),
            .I(o_One_Sec_Pulse));
    InMux I__1470 (
            .O(N__9627),
            .I(N__9624));
    LocalMux I__1469 (
            .O(N__9624),
            .I(N__9621));
    Odrv4 I__1468 (
            .O(N__9621),
            .I(\Lab_UT.bcd2segment1.m59_bmZ0 ));
    InMux I__1467 (
            .O(N__9618),
            .I(N__9615));
    LocalMux I__1466 (
            .O(N__9615),
            .I(\Lab_UT.bcd2segment1.m52_amZ0 ));
    InMux I__1465 (
            .O(N__9612),
            .I(N__9609));
    LocalMux I__1464 (
            .O(N__9609),
            .I(N__9606));
    Odrv4 I__1463 (
            .O(N__9606),
            .I(\Lab_UT.alarmcharZ0Z_0 ));
    CascadeMux I__1462 (
            .O(N__9603),
            .I(N__9600));
    InMux I__1461 (
            .O(N__9600),
            .I(N__9594));
    InMux I__1460 (
            .O(N__9599),
            .I(N__9594));
    LocalMux I__1459 (
            .O(N__9594),
            .I(N__9591));
    Span4Mux_h I__1458 (
            .O(N__9591),
            .I(N__9587));
    InMux I__1457 (
            .O(N__9590),
            .I(N__9584));
    Odrv4 I__1456 (
            .O(N__9587),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ));
    LocalMux I__1455 (
            .O(N__9584),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ));
    InMux I__1454 (
            .O(N__9579),
            .I(N__9573));
    InMux I__1453 (
            .O(N__9578),
            .I(N__9573));
    LocalMux I__1452 (
            .O(N__9573),
            .I(N__9570));
    Span4Mux_h I__1451 (
            .O(N__9570),
            .I(N__9565));
    InMux I__1450 (
            .O(N__9569),
            .I(N__9562));
    InMux I__1449 (
            .O(N__9568),
            .I(N__9559));
    Odrv4 I__1448 (
            .O(N__9565),
            .I(\Lab_UT.dictrl.next_alarmstate_1 ));
    LocalMux I__1447 (
            .O(N__9562),
            .I(\Lab_UT.dictrl.next_alarmstate_1 ));
    LocalMux I__1446 (
            .O(N__9559),
            .I(\Lab_UT.dictrl.next_alarmstate_1 ));
    CascadeMux I__1445 (
            .O(N__9552),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_ ));
    InMux I__1444 (
            .O(N__9549),
            .I(N__9546));
    LocalMux I__1443 (
            .O(N__9546),
            .I(N__9543));
    Odrv4 I__1442 (
            .O(N__9543),
            .I(\Lab_UT.bcd2segment1.m59_amZ0 ));
    InMux I__1441 (
            .O(N__9540),
            .I(N__9537));
    LocalMux I__1440 (
            .O(N__9537),
            .I(\Lab_UT.bcd2segment1.m68_bmZ0 ));
    InMux I__1439 (
            .O(N__9534),
            .I(N__9531));
    LocalMux I__1438 (
            .O(N__9531),
            .I(\uu2.un28_w_addr_user_i_0_a2Z0Z_4 ));
    InMux I__1437 (
            .O(N__9528),
            .I(N__9525));
    LocalMux I__1436 (
            .O(N__9525),
            .I(N__9520));
    InMux I__1435 (
            .O(N__9524),
            .I(N__9517));
    InMux I__1434 (
            .O(N__9523),
            .I(N__9514));
    Odrv4 I__1433 (
            .O(N__9520),
            .I(L3_tx_data_3));
    LocalMux I__1432 (
            .O(N__9517),
            .I(L3_tx_data_3));
    LocalMux I__1431 (
            .O(N__9514),
            .I(L3_tx_data_3));
    InMux I__1430 (
            .O(N__9507),
            .I(N__9503));
    CascadeMux I__1429 (
            .O(N__9506),
            .I(N__9499));
    LocalMux I__1428 (
            .O(N__9503),
            .I(N__9496));
    InMux I__1427 (
            .O(N__9502),
            .I(N__9493));
    InMux I__1426 (
            .O(N__9499),
            .I(N__9490));
    Odrv4 I__1425 (
            .O(N__9496),
            .I(L3_tx_data_4));
    LocalMux I__1424 (
            .O(N__9493),
            .I(L3_tx_data_4));
    LocalMux I__1423 (
            .O(N__9490),
            .I(L3_tx_data_4));
    InMux I__1422 (
            .O(N__9483),
            .I(N__9478));
    InMux I__1421 (
            .O(N__9482),
            .I(N__9475));
    InMux I__1420 (
            .O(N__9481),
            .I(N__9472));
    LocalMux I__1419 (
            .O(N__9478),
            .I(L3_tx_data_0));
    LocalMux I__1418 (
            .O(N__9475),
            .I(L3_tx_data_0));
    LocalMux I__1417 (
            .O(N__9472),
            .I(L3_tx_data_0));
    CascadeMux I__1416 (
            .O(N__9465),
            .I(\uu2.w_data_i_o2_4Z0Z_0_cascade_ ));
    CascadeMux I__1415 (
            .O(N__9462),
            .I(N_96_cascade_));
    CascadeMux I__1414 (
            .O(N__9459),
            .I(\uu2.un21_w_addr_displaying_i_cascade_ ));
    CascadeMux I__1413 (
            .O(N__9456),
            .I(N__9453));
    InMux I__1412 (
            .O(N__9453),
            .I(N__9450));
    LocalMux I__1411 (
            .O(N__9450),
            .I(N__9447));
    Span4Mux_v I__1410 (
            .O(N__9447),
            .I(N__9444));
    Odrv4 I__1409 (
            .O(N__9444),
            .I(\Lab_UT.alarmcharZ0Z_5 ));
    InMux I__1408 (
            .O(N__9441),
            .I(N__9438));
    LocalMux I__1407 (
            .O(N__9438),
            .I(\uu2.mem0.N_13_1_0_0 ));
    CascadeMux I__1406 (
            .O(N__9435),
            .I(\uu2.mem0.i14_mux_0_0_0_cascade_ ));
    InMux I__1405 (
            .O(N__9432),
            .I(N__9429));
    LocalMux I__1404 (
            .O(N__9429),
            .I(\uu2.mem0.N_8_0_0_1 ));
    CascadeMux I__1403 (
            .O(N__9426),
            .I(N__9423));
    InMux I__1402 (
            .O(N__9423),
            .I(N__9420));
    LocalMux I__1401 (
            .O(N__9420),
            .I(\Lab_UT.alarmcharZ0Z_6 ));
    CascadeMux I__1400 (
            .O(N__9417),
            .I(N__9413));
    CascadeMux I__1399 (
            .O(N__9416),
            .I(N__9410));
    InMux I__1398 (
            .O(N__9413),
            .I(N__9405));
    InMux I__1397 (
            .O(N__9410),
            .I(N__9405));
    LocalMux I__1396 (
            .O(N__9405),
            .I(N__9401));
    InMux I__1395 (
            .O(N__9404),
            .I(N__9398));
    Odrv4 I__1394 (
            .O(N__9401),
            .I(\uu2.N_155 ));
    LocalMux I__1393 (
            .O(N__9398),
            .I(\uu2.N_155 ));
    InMux I__1392 (
            .O(N__9393),
            .I(N__9386));
    InMux I__1391 (
            .O(N__9392),
            .I(N__9386));
    InMux I__1390 (
            .O(N__9391),
            .I(N__9383));
    LocalMux I__1389 (
            .O(N__9386),
            .I(\uu2.N_106 ));
    LocalMux I__1388 (
            .O(N__9383),
            .I(\uu2.N_106 ));
    CascadeMux I__1387 (
            .O(N__9378),
            .I(N__9373));
    InMux I__1386 (
            .O(N__9377),
            .I(N__9369));
    InMux I__1385 (
            .O(N__9376),
            .I(N__9366));
    InMux I__1384 (
            .O(N__9373),
            .I(N__9361));
    InMux I__1383 (
            .O(N__9372),
            .I(N__9361));
    LocalMux I__1382 (
            .O(N__9369),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1381 (
            .O(N__9366),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1380 (
            .O(N__9361),
            .I(\uu2.w_addr_userZ0Z_7 ));
    CascadeMux I__1379 (
            .O(N__9354),
            .I(N__9351));
    InMux I__1378 (
            .O(N__9351),
            .I(N__9348));
    LocalMux I__1377 (
            .O(N__9348),
            .I(N__9343));
    InMux I__1376 (
            .O(N__9347),
            .I(N__9340));
    InMux I__1375 (
            .O(N__9346),
            .I(N__9337));
    Odrv12 I__1374 (
            .O(N__9343),
            .I(\uu2.N_102 ));
    LocalMux I__1373 (
            .O(N__9340),
            .I(\uu2.N_102 ));
    LocalMux I__1372 (
            .O(N__9337),
            .I(\uu2.N_102 ));
    CascadeMux I__1371 (
            .O(N__9330),
            .I(N__9326));
    CascadeMux I__1370 (
            .O(N__9329),
            .I(N__9321));
    InMux I__1369 (
            .O(N__9326),
            .I(N__9317));
    InMux I__1368 (
            .O(N__9325),
            .I(N__9312));
    InMux I__1367 (
            .O(N__9324),
            .I(N__9312));
    InMux I__1366 (
            .O(N__9321),
            .I(N__9309));
    InMux I__1365 (
            .O(N__9320),
            .I(N__9305));
    LocalMux I__1364 (
            .O(N__9317),
            .I(N__9302));
    LocalMux I__1363 (
            .O(N__9312),
            .I(N__9297));
    LocalMux I__1362 (
            .O(N__9309),
            .I(N__9297));
    InMux I__1361 (
            .O(N__9308),
            .I(N__9294));
    LocalMux I__1360 (
            .O(N__9305),
            .I(\uu2.w_addr_userZ0Z_3 ));
    Odrv4 I__1359 (
            .O(N__9302),
            .I(\uu2.w_addr_userZ0Z_3 ));
    Odrv12 I__1358 (
            .O(N__9297),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1357 (
            .O(N__9294),
            .I(\uu2.w_addr_userZ0Z_3 ));
    InMux I__1356 (
            .O(N__9285),
            .I(N__9276));
    InMux I__1355 (
            .O(N__9284),
            .I(N__9265));
    InMux I__1354 (
            .O(N__9283),
            .I(N__9265));
    InMux I__1353 (
            .O(N__9282),
            .I(N__9265));
    InMux I__1352 (
            .O(N__9281),
            .I(N__9265));
    InMux I__1351 (
            .O(N__9280),
            .I(N__9265));
    CascadeMux I__1350 (
            .O(N__9279),
            .I(N__9262));
    LocalMux I__1349 (
            .O(N__9276),
            .I(N__9254));
    LocalMux I__1348 (
            .O(N__9265),
            .I(N__9254));
    InMux I__1347 (
            .O(N__9262),
            .I(N__9245));
    InMux I__1346 (
            .O(N__9261),
            .I(N__9245));
    InMux I__1345 (
            .O(N__9260),
            .I(N__9245));
    InMux I__1344 (
            .O(N__9259),
            .I(N__9245));
    Odrv4 I__1343 (
            .O(N__9254),
            .I(\uu2.N_97 ));
    LocalMux I__1342 (
            .O(N__9245),
            .I(\uu2.N_97 ));
    CascadeMux I__1341 (
            .O(N__9240),
            .I(N__9237));
    InMux I__1340 (
            .O(N__9237),
            .I(N__9228));
    InMux I__1339 (
            .O(N__9236),
            .I(N__9228));
    InMux I__1338 (
            .O(N__9235),
            .I(N__9225));
    InMux I__1337 (
            .O(N__9234),
            .I(N__9222));
    InMux I__1336 (
            .O(N__9233),
            .I(N__9219));
    LocalMux I__1335 (
            .O(N__9228),
            .I(N__9216));
    LocalMux I__1334 (
            .O(N__9225),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__1333 (
            .O(N__9222),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__1332 (
            .O(N__9219),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__1331 (
            .O(N__9216),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CEMux I__1330 (
            .O(N__9207),
            .I(N__9204));
    LocalMux I__1329 (
            .O(N__9204),
            .I(N__9201));
    Span4Mux_v I__1328 (
            .O(N__9201),
            .I(N__9198));
    Span4Mux_s2_v I__1327 (
            .O(N__9198),
            .I(N__9195));
    Odrv4 I__1326 (
            .O(N__9195),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    InMux I__1325 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__1324 (
            .O(N__9189),
            .I(N__9186));
    Odrv4 I__1323 (
            .O(N__9186),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_12 ));
    CascadeMux I__1322 (
            .O(N__9183),
            .I(\uu2.N_41_0_cascade_ ));
    InMux I__1321 (
            .O(N__9180),
            .I(N__9177));
    LocalMux I__1320 (
            .O(N__9177),
            .I(\uu2.N_132_mux ));
    CascadeMux I__1319 (
            .O(N__9174),
            .I(\uu2.N_132_mux_cascade_ ));
    InMux I__1318 (
            .O(N__9171),
            .I(N__9168));
    LocalMux I__1317 (
            .O(N__9168),
            .I(N__9165));
    Span4Mux_h I__1316 (
            .O(N__9165),
            .I(N__9162));
    Odrv4 I__1315 (
            .O(N__9162),
            .I(\uu2.mem0.N_94_i ));
    CascadeMux I__1314 (
            .O(N__9159),
            .I(N__9156));
    InMux I__1313 (
            .O(N__9156),
            .I(N__9153));
    LocalMux I__1312 (
            .O(N__9153),
            .I(N__9149));
    InMux I__1311 (
            .O(N__9152),
            .I(N__9146));
    Span4Mux_v I__1310 (
            .O(N__9149),
            .I(N__9143));
    LocalMux I__1309 (
            .O(N__9146),
            .I(\uu2.N_15_i ));
    Odrv4 I__1308 (
            .O(N__9143),
            .I(\uu2.N_15_i ));
    InMux I__1307 (
            .O(N__9138),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__1306 (
            .O(N__9135),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__1305 (
            .O(N__9132),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__1304 (
            .O(N__9129),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__1303 (
            .O(N__9126),
            .I(N__9123));
    InMux I__1302 (
            .O(N__9123),
            .I(N__9117));
    InMux I__1301 (
            .O(N__9122),
            .I(N__9117));
    LocalMux I__1300 (
            .O(N__9117),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1299 (
            .O(N__9114),
            .I(N__9111));
    InMux I__1298 (
            .O(N__9111),
            .I(N__9105));
    InMux I__1297 (
            .O(N__9110),
            .I(N__9105));
    LocalMux I__1296 (
            .O(N__9105),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1295 (
            .O(N__9102),
            .I(N__9098));
    InMux I__1294 (
            .O(N__9101),
            .I(N__9095));
    InMux I__1293 (
            .O(N__9098),
            .I(N__9092));
    LocalMux I__1292 (
            .O(N__9095),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__1291 (
            .O(N__9092),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__1290 (
            .O(N__9087),
            .I(N__9084));
    InMux I__1289 (
            .O(N__9084),
            .I(N__9078));
    InMux I__1288 (
            .O(N__9083),
            .I(N__9078));
    LocalMux I__1287 (
            .O(N__9078),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1286 (
            .O(N__9075),
            .I(N__9069));
    InMux I__1285 (
            .O(N__9074),
            .I(N__9069));
    LocalMux I__1284 (
            .O(N__9069),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1283 (
            .O(N__9066),
            .I(N__9058));
    InMux I__1282 (
            .O(N__9065),
            .I(N__9058));
    InMux I__1281 (
            .O(N__9064),
            .I(N__9055));
    InMux I__1280 (
            .O(N__9063),
            .I(N__9052));
    LocalMux I__1279 (
            .O(N__9058),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1278 (
            .O(N__9055),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1277 (
            .O(N__9052),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1276 (
            .O(N__9045),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ));
    CascadeMux I__1275 (
            .O(N__9042),
            .I(N__9038));
    InMux I__1274 (
            .O(N__9041),
            .I(N__9034));
    InMux I__1273 (
            .O(N__9038),
            .I(N__9029));
    InMux I__1272 (
            .O(N__9037),
            .I(N__9029));
    LocalMux I__1271 (
            .O(N__9034),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1270 (
            .O(N__9029),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1269 (
            .O(N__9024),
            .I(N__9018));
    InMux I__1268 (
            .O(N__9023),
            .I(N__9011));
    InMux I__1267 (
            .O(N__9022),
            .I(N__9011));
    InMux I__1266 (
            .O(N__9021),
            .I(N__9011));
    LocalMux I__1265 (
            .O(N__9018),
            .I(N__9008));
    LocalMux I__1264 (
            .O(N__9011),
            .I(\buart.Z_tx.ser_clk ));
    Odrv4 I__1263 (
            .O(N__9008),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__1262 (
            .O(N__9003),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    CascadeMux I__1261 (
            .O(N__9000),
            .I(N__8995));
    CascadeMux I__1260 (
            .O(N__8999),
            .I(N__8992));
    CascadeMux I__1259 (
            .O(N__8998),
            .I(N__8989));
    InMux I__1258 (
            .O(N__8995),
            .I(N__8982));
    InMux I__1257 (
            .O(N__8992),
            .I(N__8982));
    InMux I__1256 (
            .O(N__8989),
            .I(N__8982));
    LocalMux I__1255 (
            .O(N__8982),
            .I(\uu2.l_countZ0Z_9 ));
    CascadeMux I__1254 (
            .O(N__8979),
            .I(N__8975));
    InMux I__1253 (
            .O(N__8978),
            .I(N__8971));
    InMux I__1252 (
            .O(N__8975),
            .I(N__8966));
    InMux I__1251 (
            .O(N__8974),
            .I(N__8966));
    LocalMux I__1250 (
            .O(N__8971),
            .I(N__8963));
    LocalMux I__1249 (
            .O(N__8966),
            .I(\uu2.l_countZ0Z_7 ));
    Odrv4 I__1248 (
            .O(N__8963),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__1247 (
            .O(N__8958),
            .I(N__8952));
    InMux I__1246 (
            .O(N__8957),
            .I(N__8952));
    LocalMux I__1245 (
            .O(N__8952),
            .I(\uu2.un1_l_count_1_3 ));
    InMux I__1244 (
            .O(N__8949),
            .I(N__8940));
    InMux I__1243 (
            .O(N__8948),
            .I(N__8940));
    InMux I__1242 (
            .O(N__8947),
            .I(N__8937));
    InMux I__1241 (
            .O(N__8946),
            .I(N__8932));
    InMux I__1240 (
            .O(N__8945),
            .I(N__8932));
    LocalMux I__1239 (
            .O(N__8940),
            .I(N__8929));
    LocalMux I__1238 (
            .O(N__8937),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1237 (
            .O(N__8932),
            .I(\uu2.l_countZ0Z_1 ));
    Odrv4 I__1236 (
            .O(N__8929),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__1235 (
            .O(N__8922),
            .I(N__8914));
    InMux I__1234 (
            .O(N__8921),
            .I(N__8914));
    InMux I__1233 (
            .O(N__8920),
            .I(N__8907));
    InMux I__1232 (
            .O(N__8919),
            .I(N__8907));
    LocalMux I__1231 (
            .O(N__8914),
            .I(N__8904));
    InMux I__1230 (
            .O(N__8913),
            .I(N__8899));
    InMux I__1229 (
            .O(N__8912),
            .I(N__8899));
    LocalMux I__1228 (
            .O(N__8907),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__1227 (
            .O(N__8904),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1226 (
            .O(N__8899),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__1225 (
            .O(N__8892),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__1224 (
            .O(N__8889),
            .I(N__8878));
    CascadeMux I__1223 (
            .O(N__8888),
            .I(N__8875));
    InMux I__1222 (
            .O(N__8887),
            .I(N__8853));
    InMux I__1221 (
            .O(N__8886),
            .I(N__8853));
    InMux I__1220 (
            .O(N__8885),
            .I(N__8853));
    InMux I__1219 (
            .O(N__8884),
            .I(N__8853));
    InMux I__1218 (
            .O(N__8883),
            .I(N__8853));
    InMux I__1217 (
            .O(N__8882),
            .I(N__8853));
    InMux I__1216 (
            .O(N__8881),
            .I(N__8853));
    LocalMux I__1215 (
            .O(N__8878),
            .I(N__8850));
    InMux I__1214 (
            .O(N__8875),
            .I(N__8845));
    InMux I__1213 (
            .O(N__8874),
            .I(N__8845));
    InMux I__1212 (
            .O(N__8873),
            .I(N__8838));
    InMux I__1211 (
            .O(N__8872),
            .I(N__8838));
    InMux I__1210 (
            .O(N__8871),
            .I(N__8838));
    InMux I__1209 (
            .O(N__8870),
            .I(N__8835));
    InMux I__1208 (
            .O(N__8869),
            .I(N__8832));
    CascadeMux I__1207 (
            .O(N__8868),
            .I(N__8829));
    LocalMux I__1206 (
            .O(N__8853),
            .I(N__8826));
    Span4Mux_s2_h I__1205 (
            .O(N__8850),
            .I(N__8821));
    LocalMux I__1204 (
            .O(N__8845),
            .I(N__8821));
    LocalMux I__1203 (
            .O(N__8838),
            .I(N__8818));
    LocalMux I__1202 (
            .O(N__8835),
            .I(N__8813));
    LocalMux I__1201 (
            .O(N__8832),
            .I(N__8813));
    InMux I__1200 (
            .O(N__8829),
            .I(N__8810));
    Span4Mux_s3_h I__1199 (
            .O(N__8826),
            .I(N__8807));
    Span4Mux_v I__1198 (
            .O(N__8821),
            .I(N__8804));
    Span4Mux_s3_h I__1197 (
            .O(N__8818),
            .I(N__8801));
    Span4Mux_h I__1196 (
            .O(N__8813),
            .I(N__8798));
    LocalMux I__1195 (
            .O(N__8810),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1194 (
            .O(N__8807),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1193 (
            .O(N__8804),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1192 (
            .O(N__8801),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1191 (
            .O(N__8798),
            .I(vbuf_tx_data_rdy));
    InMux I__1190 (
            .O(N__8787),
            .I(N__8783));
    CascadeMux I__1189 (
            .O(N__8786),
            .I(N__8780));
    LocalMux I__1188 (
            .O(N__8783),
            .I(N__8775));
    InMux I__1187 (
            .O(N__8780),
            .I(N__8770));
    InMux I__1186 (
            .O(N__8779),
            .I(N__8770));
    InMux I__1185 (
            .O(N__8778),
            .I(N__8767));
    Odrv4 I__1184 (
            .O(N__8775),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__1183 (
            .O(N__8770),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__1182 (
            .O(N__8767),
            .I(\uu0.l_countZ0Z_10 ));
    InMux I__1181 (
            .O(N__8760),
            .I(N__8757));
    LocalMux I__1180 (
            .O(N__8757),
            .I(N__8751));
    InMux I__1179 (
            .O(N__8756),
            .I(N__8746));
    InMux I__1178 (
            .O(N__8755),
            .I(N__8743));
    InMux I__1177 (
            .O(N__8754),
            .I(N__8740));
    Span4Mux_h I__1176 (
            .O(N__8751),
            .I(N__8737));
    InMux I__1175 (
            .O(N__8750),
            .I(N__8732));
    InMux I__1174 (
            .O(N__8749),
            .I(N__8732));
    LocalMux I__1173 (
            .O(N__8746),
            .I(N__8727));
    LocalMux I__1172 (
            .O(N__8743),
            .I(N__8727));
    LocalMux I__1171 (
            .O(N__8740),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1170 (
            .O(N__8737),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1169 (
            .O(N__8732),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1168 (
            .O(N__8727),
            .I(\uu0.l_countZ0Z_8 ));
    InMux I__1167 (
            .O(N__8718),
            .I(N__8715));
    LocalMux I__1166 (
            .O(N__8715),
            .I(N__8711));
    InMux I__1165 (
            .O(N__8714),
            .I(N__8705));
    Span4Mux_h I__1164 (
            .O(N__8711),
            .I(N__8702));
    InMux I__1163 (
            .O(N__8710),
            .I(N__8697));
    InMux I__1162 (
            .O(N__8709),
            .I(N__8697));
    InMux I__1161 (
            .O(N__8708),
            .I(N__8694));
    LocalMux I__1160 (
            .O(N__8705),
            .I(\uu0.l_countZ0Z_9 ));
    Odrv4 I__1159 (
            .O(N__8702),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1158 (
            .O(N__8697),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1157 (
            .O(N__8694),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__1156 (
            .O(N__8685),
            .I(N__8682));
    LocalMux I__1155 (
            .O(N__8682),
            .I(N__8679));
    Span4Mux_s3_h I__1154 (
            .O(N__8679),
            .I(N__8676));
    Odrv4 I__1153 (
            .O(N__8676),
            .I(\uu0.un143_ci_0 ));
    CascadeMux I__1152 (
            .O(N__8673),
            .I(\uu2.un1_l_count_1_2_0_cascade_ ));
    InMux I__1151 (
            .O(N__8670),
            .I(N__8666));
    InMux I__1150 (
            .O(N__8669),
            .I(N__8663));
    LocalMux I__1149 (
            .O(N__8666),
            .I(N__8660));
    LocalMux I__1148 (
            .O(N__8663),
            .I(N__8655));
    Span4Mux_s3_h I__1147 (
            .O(N__8660),
            .I(N__8655));
    Odrv4 I__1146 (
            .O(N__8655),
            .I(\uu2.un1_l_count_1_0 ));
    CascadeMux I__1145 (
            .O(N__8652),
            .I(\uu2.un1_l_count_2_2_cascade_ ));
    CascadeMux I__1144 (
            .O(N__8649),
            .I(\resetGen.reset_count_2_0_4_cascade_ ));
    InMux I__1143 (
            .O(N__8646),
            .I(N__8643));
    LocalMux I__1142 (
            .O(N__8643),
            .I(N__8640));
    Odrv4 I__1141 (
            .O(N__8640),
            .I(\Lab_UT.alarmchar10 ));
    CascadeMux I__1140 (
            .O(N__8637),
            .I(N__8634));
    InMux I__1139 (
            .O(N__8634),
            .I(N__8631));
    LocalMux I__1138 (
            .O(N__8631),
            .I(\Lab_UT.alarmcharZ0Z_4 ));
    CascadeMux I__1137 (
            .O(N__8628),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__1136 (
            .O(N__8625),
            .I(N__8621));
    InMux I__1135 (
            .O(N__8624),
            .I(N__8618));
    LocalMux I__1134 (
            .O(N__8621),
            .I(\resetGen.reset_countZ0Z_3 ));
    LocalMux I__1133 (
            .O(N__8618),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__1132 (
            .O(N__8613),
            .I(N__8606));
    InMux I__1131 (
            .O(N__8612),
            .I(N__8606));
    InMux I__1130 (
            .O(N__8611),
            .I(N__8603));
    LocalMux I__1129 (
            .O(N__8606),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__1128 (
            .O(N__8603),
            .I(\resetGen.reset_countZ0Z_1 ));
    InMux I__1127 (
            .O(N__8598),
            .I(N__8595));
    LocalMux I__1126 (
            .O(N__8595),
            .I(\resetGen.un241_ci ));
    CascadeMux I__1125 (
            .O(N__8592),
            .I(\resetGen.un241_ci_cascade_ ));
    InMux I__1124 (
            .O(N__8589),
            .I(N__8584));
    InMux I__1123 (
            .O(N__8588),
            .I(N__8581));
    InMux I__1122 (
            .O(N__8587),
            .I(N__8578));
    LocalMux I__1121 (
            .O(N__8584),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1120 (
            .O(N__8581),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1119 (
            .O(N__8578),
            .I(\resetGen.reset_countZ0Z_2 ));
    CascadeMux I__1118 (
            .O(N__8571),
            .I(N__8568));
    InMux I__1117 (
            .O(N__8568),
            .I(N__8556));
    InMux I__1116 (
            .O(N__8567),
            .I(N__8556));
    InMux I__1115 (
            .O(N__8566),
            .I(N__8556));
    InMux I__1114 (
            .O(N__8565),
            .I(N__8556));
    LocalMux I__1113 (
            .O(N__8556),
            .I(\resetGen.reset_countZ0Z_0 ));
    CascadeMux I__1112 (
            .O(N__8553),
            .I(\uu2.un28_w_addr_user_i_0_cascade_ ));
    InMux I__1111 (
            .O(N__8550),
            .I(N__8547));
    LocalMux I__1110 (
            .O(N__8547),
            .I(N__8541));
    InMux I__1109 (
            .O(N__8546),
            .I(N__8536));
    InMux I__1108 (
            .O(N__8545),
            .I(N__8536));
    InMux I__1107 (
            .O(N__8544),
            .I(N__8533));
    Odrv4 I__1106 (
            .O(N__8541),
            .I(\uu2.un28_w_addr_user_i_0 ));
    LocalMux I__1105 (
            .O(N__8536),
            .I(\uu2.un28_w_addr_user_i_0 ));
    LocalMux I__1104 (
            .O(N__8533),
            .I(\uu2.un28_w_addr_user_i_0 ));
    InMux I__1103 (
            .O(N__8526),
            .I(N__8523));
    LocalMux I__1102 (
            .O(N__8523),
            .I(N__8520));
    Odrv4 I__1101 (
            .O(N__8520),
            .I(\uu2.N_105 ));
    CascadeMux I__1100 (
            .O(N__8517),
            .I(N__8514));
    InMux I__1099 (
            .O(N__8514),
            .I(N__8508));
    InMux I__1098 (
            .O(N__8513),
            .I(N__8503));
    InMux I__1097 (
            .O(N__8512),
            .I(N__8503));
    InMux I__1096 (
            .O(N__8511),
            .I(N__8500));
    LocalMux I__1095 (
            .O(N__8508),
            .I(N__8495));
    LocalMux I__1094 (
            .O(N__8503),
            .I(N__8495));
    LocalMux I__1093 (
            .O(N__8500),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__1092 (
            .O(N__8495),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__1091 (
            .O(N__8490),
            .I(\uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_ ));
    InMux I__1090 (
            .O(N__8487),
            .I(N__8484));
    LocalMux I__1089 (
            .O(N__8484),
            .I(N__8481));
    Odrv4 I__1088 (
            .O(N__8481),
            .I(\Lab_UT.alarmchar_2_1_1 ));
    CascadeMux I__1087 (
            .O(N__8478),
            .I(N__8475));
    InMux I__1086 (
            .O(N__8475),
            .I(N__8472));
    LocalMux I__1085 (
            .O(N__8472),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_4 ));
    InMux I__1084 (
            .O(N__8469),
            .I(N__8466));
    LocalMux I__1083 (
            .O(N__8466),
            .I(\uu2.w_addr_user_3_i_a2_3_6 ));
    CascadeMux I__1082 (
            .O(N__8463),
            .I(\uu2.mem0.g1_3_0_cascade_ ));
    InMux I__1081 (
            .O(N__8460),
            .I(N__8457));
    LocalMux I__1080 (
            .O(N__8457),
            .I(\uu2.mem0.N_63_0_i ));
    InMux I__1079 (
            .O(N__8454),
            .I(N__8451));
    LocalMux I__1078 (
            .O(N__8451),
            .I(\uu2.mem0.G_17_0_0_0 ));
    CascadeMux I__1077 (
            .O(N__8448),
            .I(N__8444));
    CascadeMux I__1076 (
            .O(N__8447),
            .I(N__8441));
    InMux I__1075 (
            .O(N__8444),
            .I(N__8436));
    InMux I__1074 (
            .O(N__8441),
            .I(N__8436));
    LocalMux I__1073 (
            .O(N__8436),
            .I(N_72_mux));
    CascadeMux I__1072 (
            .O(N__8433),
            .I(N__8430));
    InMux I__1071 (
            .O(N__8430),
            .I(N__8427));
    LocalMux I__1070 (
            .O(N__8427),
            .I(N__8424));
    Span4Mux_s3_h I__1069 (
            .O(N__8424),
            .I(N__8421));
    Odrv4 I__1068 (
            .O(N__8421),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_3 ));
    InMux I__1067 (
            .O(N__8418),
            .I(N__8415));
    LocalMux I__1066 (
            .O(N__8415),
            .I(\uu2.w_addr_user_3_i_a2_2_6 ));
    CascadeMux I__1065 (
            .O(N__8412),
            .I(N__8409));
    InMux I__1064 (
            .O(N__8409),
            .I(N__8406));
    LocalMux I__1063 (
            .O(N__8406),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_2 ));
    CascadeMux I__1062 (
            .O(N__8403),
            .I(N__8400));
    InMux I__1061 (
            .O(N__8400),
            .I(N__8397));
    LocalMux I__1060 (
            .O(N__8397),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_6 ));
    CascadeMux I__1059 (
            .O(N__8394),
            .I(N__8391));
    InMux I__1058 (
            .O(N__8391),
            .I(N__8388));
    LocalMux I__1057 (
            .O(N__8388),
            .I(N__8385));
    Odrv4 I__1056 (
            .O(N__8385),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_7 ));
    CascadeMux I__1055 (
            .O(N__8382),
            .I(\uu2.N_102_cascade_ ));
    CascadeMux I__1054 (
            .O(N__8379),
            .I(N__8376));
    InMux I__1053 (
            .O(N__8376),
            .I(N__8373));
    LocalMux I__1052 (
            .O(N__8373),
            .I(\uu2.N_61_i ));
    CascadeMux I__1051 (
            .O(N__8370),
            .I(N__8364));
    CascadeMux I__1050 (
            .O(N__8369),
            .I(N__8361));
    InMux I__1049 (
            .O(N__8368),
            .I(N__8358));
    InMux I__1048 (
            .O(N__8367),
            .I(N__8351));
    InMux I__1047 (
            .O(N__8364),
            .I(N__8351));
    InMux I__1046 (
            .O(N__8361),
            .I(N__8351));
    LocalMux I__1045 (
            .O(N__8358),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__1044 (
            .O(N__8351),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CascadeMux I__1043 (
            .O(N__8346),
            .I(\buart.Z_tx.un1_bitcount_c3_cascade_ ));
    InMux I__1042 (
            .O(N__8343),
            .I(N__8339));
    InMux I__1041 (
            .O(N__8342),
            .I(N__8336));
    LocalMux I__1040 (
            .O(N__8339),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__1039 (
            .O(N__8336),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__1038 (
            .O(N__8331),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    InMux I__1037 (
            .O(N__8328),
            .I(N__8321));
    InMux I__1036 (
            .O(N__8327),
            .I(N__8318));
    InMux I__1035 (
            .O(N__8326),
            .I(N__8311));
    InMux I__1034 (
            .O(N__8325),
            .I(N__8311));
    InMux I__1033 (
            .O(N__8324),
            .I(N__8311));
    LocalMux I__1032 (
            .O(N__8321),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__1031 (
            .O(N__8318),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__1030 (
            .O(N__8311),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    InMux I__1029 (
            .O(N__8304),
            .I(N__8292));
    InMux I__1028 (
            .O(N__8303),
            .I(N__8292));
    InMux I__1027 (
            .O(N__8302),
            .I(N__8292));
    InMux I__1026 (
            .O(N__8301),
            .I(N__8292));
    LocalMux I__1025 (
            .O(N__8292),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__1024 (
            .O(N__8289),
            .I(N__8284));
    InMux I__1023 (
            .O(N__8288),
            .I(N__8279));
    InMux I__1022 (
            .O(N__8287),
            .I(N__8274));
    InMux I__1021 (
            .O(N__8284),
            .I(N__8274));
    InMux I__1020 (
            .O(N__8283),
            .I(N__8269));
    InMux I__1019 (
            .O(N__8282),
            .I(N__8269));
    LocalMux I__1018 (
            .O(N__8279),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1017 (
            .O(N__8274),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1016 (
            .O(N__8269),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__1015 (
            .O(N__8262),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    CascadeMux I__1014 (
            .O(N__8259),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ));
    InMux I__1013 (
            .O(N__8256),
            .I(N__8247));
    InMux I__1012 (
            .O(N__8255),
            .I(N__8247));
    InMux I__1011 (
            .O(N__8254),
            .I(N__8247));
    LocalMux I__1010 (
            .O(N__8247),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    InMux I__1009 (
            .O(N__8244),
            .I(N__8241));
    LocalMux I__1008 (
            .O(N__8241),
            .I(N__8238));
    Span4Mux_h I__1007 (
            .O(N__8238),
            .I(N__8235));
    Span4Mux_v I__1006 (
            .O(N__8235),
            .I(N__8232));
    Odrv4 I__1005 (
            .O(N__8232),
            .I(\Lab_UT.alarmchar10_i_2 ));
    CascadeMux I__1004 (
            .O(N__8229),
            .I(N__8224));
    InMux I__1003 (
            .O(N__8228),
            .I(N__8219));
    InMux I__1002 (
            .O(N__8227),
            .I(N__8219));
    InMux I__1001 (
            .O(N__8224),
            .I(N__8216));
    LocalMux I__1000 (
            .O(N__8219),
            .I(\uu0.l_countZ0Z_17 ));
    LocalMux I__999 (
            .O(N__8216),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__998 (
            .O(N__8211),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__997 (
            .O(N__8208),
            .I(N__8204));
    InMux I__996 (
            .O(N__8207),
            .I(N__8201));
    LocalMux I__995 (
            .O(N__8204),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__994 (
            .O(N__8201),
            .I(\uu0.l_countZ0Z_18 ));
    CEMux I__993 (
            .O(N__8196),
            .I(N__8181));
    CEMux I__992 (
            .O(N__8195),
            .I(N__8181));
    CEMux I__991 (
            .O(N__8194),
            .I(N__8181));
    CEMux I__990 (
            .O(N__8193),
            .I(N__8181));
    CEMux I__989 (
            .O(N__8192),
            .I(N__8181));
    GlobalMux I__988 (
            .O(N__8181),
            .I(N__8178));
    gio2CtrlBuf I__987 (
            .O(N__8178),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__986 (
            .O(N__8175),
            .I(N__8170));
    InMux I__985 (
            .O(N__8174),
            .I(N__8165));
    InMux I__984 (
            .O(N__8173),
            .I(N__8165));
    InMux I__983 (
            .O(N__8170),
            .I(N__8162));
    LocalMux I__982 (
            .O(N__8165),
            .I(\uu0.l_precountZ0Z_3 ));
    LocalMux I__981 (
            .O(N__8162),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__980 (
            .O(N__8157),
            .I(N__8154));
    InMux I__979 (
            .O(N__8154),
            .I(N__8141));
    InMux I__978 (
            .O(N__8153),
            .I(N__8141));
    InMux I__977 (
            .O(N__8152),
            .I(N__8141));
    InMux I__976 (
            .O(N__8151),
            .I(N__8141));
    InMux I__975 (
            .O(N__8150),
            .I(N__8138));
    LocalMux I__974 (
            .O(N__8141),
            .I(\uu0.l_precountZ0Z_1 ));
    LocalMux I__973 (
            .O(N__8138),
            .I(\uu0.l_precountZ0Z_1 ));
    InMux I__972 (
            .O(N__8133),
            .I(N__8123));
    InMux I__971 (
            .O(N__8132),
            .I(N__8123));
    InMux I__970 (
            .O(N__8131),
            .I(N__8123));
    InMux I__969 (
            .O(N__8130),
            .I(N__8120));
    LocalMux I__968 (
            .O(N__8123),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__967 (
            .O(N__8120),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__966 (
            .O(N__8115),
            .I(N__8109));
    InMux I__965 (
            .O(N__8114),
            .I(N__8100));
    InMux I__964 (
            .O(N__8113),
            .I(N__8100));
    InMux I__963 (
            .O(N__8112),
            .I(N__8100));
    InMux I__962 (
            .O(N__8109),
            .I(N__8100));
    LocalMux I__961 (
            .O(N__8100),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__960 (
            .O(N__8097),
            .I(N__8081));
    InMux I__959 (
            .O(N__8096),
            .I(N__8081));
    InMux I__958 (
            .O(N__8095),
            .I(N__8081));
    InMux I__957 (
            .O(N__8094),
            .I(N__8081));
    InMux I__956 (
            .O(N__8093),
            .I(N__8081));
    InMux I__955 (
            .O(N__8092),
            .I(N__8078));
    LocalMux I__954 (
            .O(N__8081),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__953 (
            .O(N__8078),
            .I(\uu0.l_countZ0Z_0 ));
    CascadeMux I__952 (
            .O(N__8073),
            .I(N__8070));
    InMux I__951 (
            .O(N__8070),
            .I(N__8062));
    InMux I__950 (
            .O(N__8069),
            .I(N__8062));
    InMux I__949 (
            .O(N__8068),
            .I(N__8059));
    InMux I__948 (
            .O(N__8067),
            .I(N__8056));
    LocalMux I__947 (
            .O(N__8062),
            .I(N__8051));
    LocalMux I__946 (
            .O(N__8059),
            .I(N__8051));
    LocalMux I__945 (
            .O(N__8056),
            .I(\uu0.l_countZ0Z_16 ));
    Odrv4 I__944 (
            .O(N__8051),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__943 (
            .O(N__8046),
            .I(\uu0.un4_l_count_14_cascade_ ));
    InMux I__942 (
            .O(N__8043),
            .I(N__8033));
    InMux I__941 (
            .O(N__8042),
            .I(N__8033));
    InMux I__940 (
            .O(N__8041),
            .I(N__8033));
    InMux I__939 (
            .O(N__8040),
            .I(N__8030));
    LocalMux I__938 (
            .O(N__8033),
            .I(N__8027));
    LocalMux I__937 (
            .O(N__8030),
            .I(N__8024));
    Odrv4 I__936 (
            .O(N__8027),
            .I(\uu0.un4_l_count_0_8 ));
    Odrv12 I__935 (
            .O(N__8024),
            .I(\uu0.un4_l_count_0_8 ));
    InMux I__934 (
            .O(N__8019),
            .I(N__8016));
    LocalMux I__933 (
            .O(N__8016),
            .I(\uu0.un4_l_count_18 ));
    CascadeMux I__932 (
            .O(N__8013),
            .I(N__8006));
    InMux I__931 (
            .O(N__8012),
            .I(N__7992));
    InMux I__930 (
            .O(N__8011),
            .I(N__7992));
    InMux I__929 (
            .O(N__8010),
            .I(N__7992));
    InMux I__928 (
            .O(N__8009),
            .I(N__7992));
    InMux I__927 (
            .O(N__8006),
            .I(N__7992));
    InMux I__926 (
            .O(N__8005),
            .I(N__7992));
    LocalMux I__925 (
            .O(N__7992),
            .I(\uu0.l_precountZ0Z_0 ));
    InMux I__924 (
            .O(N__7989),
            .I(N__7985));
    InMux I__923 (
            .O(N__7988),
            .I(N__7982));
    LocalMux I__922 (
            .O(N__7985),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    LocalMux I__921 (
            .O(N__7982),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    InMux I__920 (
            .O(N__7977),
            .I(N__7974));
    LocalMux I__919 (
            .O(N__7974),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__918 (
            .O(N__7971),
            .I(N__7967));
    InMux I__917 (
            .O(N__7970),
            .I(N__7964));
    LocalMux I__916 (
            .O(N__7967),
            .I(N__7961));
    LocalMux I__915 (
            .O(N__7964),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__914 (
            .O(N__7961),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__913 (
            .O(N__7956),
            .I(N__7953));
    LocalMux I__912 (
            .O(N__7953),
            .I(N__7950));
    Odrv4 I__911 (
            .O(N__7950),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__910 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__909 (
            .O(N__7944),
            .I(\uu0.un55_ci ));
    InMux I__908 (
            .O(N__7941),
            .I(N__7936));
    InMux I__907 (
            .O(N__7940),
            .I(N__7933));
    InMux I__906 (
            .O(N__7939),
            .I(N__7930));
    LocalMux I__905 (
            .O(N__7936),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__904 (
            .O(N__7933),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__903 (
            .O(N__7930),
            .I(\uu0.l_countZ0Z_3 ));
    CascadeMux I__902 (
            .O(N__7923),
            .I(N__7919));
    CascadeMux I__901 (
            .O(N__7922),
            .I(N__7916));
    InMux I__900 (
            .O(N__7919),
            .I(N__7912));
    InMux I__899 (
            .O(N__7916),
            .I(N__7909));
    InMux I__898 (
            .O(N__7915),
            .I(N__7906));
    LocalMux I__897 (
            .O(N__7912),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__896 (
            .O(N__7909),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__895 (
            .O(N__7906),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__894 (
            .O(N__7899),
            .I(N__7891));
    InMux I__893 (
            .O(N__7898),
            .I(N__7881));
    InMux I__892 (
            .O(N__7897),
            .I(N__7881));
    InMux I__891 (
            .O(N__7896),
            .I(N__7876));
    InMux I__890 (
            .O(N__7895),
            .I(N__7876));
    InMux I__889 (
            .O(N__7894),
            .I(N__7871));
    InMux I__888 (
            .O(N__7891),
            .I(N__7871));
    InMux I__887 (
            .O(N__7890),
            .I(N__7868));
    InMux I__886 (
            .O(N__7889),
            .I(N__7859));
    InMux I__885 (
            .O(N__7888),
            .I(N__7859));
    InMux I__884 (
            .O(N__7887),
            .I(N__7859));
    InMux I__883 (
            .O(N__7886),
            .I(N__7859));
    LocalMux I__882 (
            .O(N__7881),
            .I(N__7854));
    LocalMux I__881 (
            .O(N__7876),
            .I(N__7854));
    LocalMux I__880 (
            .O(N__7871),
            .I(\uu0.un110_ci ));
    LocalMux I__879 (
            .O(N__7868),
            .I(\uu0.un110_ci ));
    LocalMux I__878 (
            .O(N__7859),
            .I(\uu0.un110_ci ));
    Odrv12 I__877 (
            .O(N__7854),
            .I(\uu0.un110_ci ));
    CascadeMux I__876 (
            .O(N__7845),
            .I(N__7841));
    CascadeMux I__875 (
            .O(N__7844),
            .I(N__7837));
    InMux I__874 (
            .O(N__7841),
            .I(N__7834));
    InMux I__873 (
            .O(N__7840),
            .I(N__7829));
    InMux I__872 (
            .O(N__7837),
            .I(N__7829));
    LocalMux I__871 (
            .O(N__7834),
            .I(\uu0.un198_ci_2 ));
    LocalMux I__870 (
            .O(N__7829),
            .I(\uu0.un198_ci_2 ));
    InMux I__869 (
            .O(N__7824),
            .I(N__7820));
    InMux I__868 (
            .O(N__7823),
            .I(N__7817));
    LocalMux I__867 (
            .O(N__7820),
            .I(\uu0.l_countZ0Z_13 ));
    LocalMux I__866 (
            .O(N__7817),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__865 (
            .O(N__7812),
            .I(N__7807));
    InMux I__864 (
            .O(N__7811),
            .I(N__7802));
    InMux I__863 (
            .O(N__7810),
            .I(N__7802));
    LocalMux I__862 (
            .O(N__7807),
            .I(\uu0.l_countZ0Z_12 ));
    LocalMux I__861 (
            .O(N__7802),
            .I(\uu0.l_countZ0Z_12 ));
    CascadeMux I__860 (
            .O(N__7797),
            .I(N__7794));
    InMux I__859 (
            .O(N__7794),
            .I(N__7790));
    InMux I__858 (
            .O(N__7793),
            .I(N__7785));
    LocalMux I__857 (
            .O(N__7790),
            .I(N__7782));
    InMux I__856 (
            .O(N__7789),
            .I(N__7777));
    InMux I__855 (
            .O(N__7788),
            .I(N__7777));
    LocalMux I__854 (
            .O(N__7785),
            .I(N__7774));
    Odrv12 I__853 (
            .O(N__7782),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__852 (
            .O(N__7777),
            .I(\uu0.un154_ci_9 ));
    Odrv4 I__851 (
            .O(N__7774),
            .I(\uu0.un154_ci_9 ));
    CascadeMux I__850 (
            .O(N__7767),
            .I(N__7764));
    InMux I__849 (
            .O(N__7764),
            .I(N__7761));
    LocalMux I__848 (
            .O(N__7761),
            .I(\uu0.un165_ci_0 ));
    InMux I__847 (
            .O(N__7758),
            .I(N__7755));
    LocalMux I__846 (
            .O(N__7755),
            .I(N__7752));
    Span4Mux_h I__845 (
            .O(N__7752),
            .I(N__7749));
    Odrv4 I__844 (
            .O(N__7749),
            .I(\uu0.sec_clkDZ0 ));
    CascadeMux I__843 (
            .O(N__7746),
            .I(N__7743));
    InMux I__842 (
            .O(N__7743),
            .I(N__7738));
    InMux I__841 (
            .O(N__7742),
            .I(N__7732));
    InMux I__840 (
            .O(N__7741),
            .I(N__7732));
    LocalMux I__839 (
            .O(N__7738),
            .I(N__7729));
    InMux I__838 (
            .O(N__7737),
            .I(N__7726));
    LocalMux I__837 (
            .O(N__7732),
            .I(N__7723));
    Odrv4 I__836 (
            .O(N__7729),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__835 (
            .O(N__7726),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__834 (
            .O(N__7723),
            .I(\uu2.r_addrZ0Z_5 ));
    CascadeMux I__833 (
            .O(N__7716),
            .I(N__7711));
    InMux I__832 (
            .O(N__7715),
            .I(N__7705));
    InMux I__831 (
            .O(N__7714),
            .I(N__7705));
    InMux I__830 (
            .O(N__7711),
            .I(N__7700));
    InMux I__829 (
            .O(N__7710),
            .I(N__7700));
    LocalMux I__828 (
            .O(N__7705),
            .I(N__7697));
    LocalMux I__827 (
            .O(N__7700),
            .I(N__7694));
    Odrv4 I__826 (
            .O(N__7697),
            .I(\uu2.un404_ci ));
    Odrv4 I__825 (
            .O(N__7694),
            .I(\uu2.un404_ci ));
    CascadeMux I__824 (
            .O(N__7689),
            .I(N__7686));
    InMux I__823 (
            .O(N__7686),
            .I(N__7679));
    InMux I__822 (
            .O(N__7685),
            .I(N__7674));
    InMux I__821 (
            .O(N__7684),
            .I(N__7674));
    InMux I__820 (
            .O(N__7683),
            .I(N__7669));
    InMux I__819 (
            .O(N__7682),
            .I(N__7669));
    LocalMux I__818 (
            .O(N__7679),
            .I(N__7664));
    LocalMux I__817 (
            .O(N__7674),
            .I(N__7664));
    LocalMux I__816 (
            .O(N__7669),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__815 (
            .O(N__7664),
            .I(\uu2.r_addrZ0Z_4 ));
    CEMux I__814 (
            .O(N__7659),
            .I(N__7656));
    LocalMux I__813 (
            .O(N__7656),
            .I(N__7652));
    CEMux I__812 (
            .O(N__7655),
            .I(N__7649));
    Span4Mux_h I__811 (
            .O(N__7652),
            .I(N__7644));
    LocalMux I__810 (
            .O(N__7649),
            .I(N__7644));
    Sp12to4 I__809 (
            .O(N__7644),
            .I(N__7641));
    Odrv12 I__808 (
            .O(N__7641),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__807 (
            .O(N__7638),
            .I(N__7635));
    InMux I__806 (
            .O(N__7635),
            .I(N__7631));
    CascadeMux I__805 (
            .O(N__7634),
            .I(N__7627));
    LocalMux I__804 (
            .O(N__7631),
            .I(N__7624));
    CascadeMux I__803 (
            .O(N__7630),
            .I(N__7621));
    InMux I__802 (
            .O(N__7627),
            .I(N__7618));
    Span4Mux_h I__801 (
            .O(N__7624),
            .I(N__7615));
    InMux I__800 (
            .O(N__7621),
            .I(N__7612));
    LocalMux I__799 (
            .O(N__7618),
            .I(N__7609));
    Odrv4 I__798 (
            .O(N__7615),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__797 (
            .O(N__7612),
            .I(\uu2.r_addrZ0Z_3 ));
    Odrv4 I__796 (
            .O(N__7609),
            .I(\uu2.r_addrZ0Z_3 ));
    CascadeMux I__795 (
            .O(N__7602),
            .I(\uu2.un404_ci_cascade_ ));
    CascadeMux I__794 (
            .O(N__7599),
            .I(N__7596));
    InMux I__793 (
            .O(N__7596),
            .I(N__7592));
    InMux I__792 (
            .O(N__7595),
            .I(N__7588));
    LocalMux I__791 (
            .O(N__7592),
            .I(N__7585));
    InMux I__790 (
            .O(N__7591),
            .I(N__7582));
    LocalMux I__789 (
            .O(N__7588),
            .I(N__7579));
    Odrv4 I__788 (
            .O(N__7585),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__787 (
            .O(N__7582),
            .I(\uu2.r_addrZ0Z_7 ));
    Odrv4 I__786 (
            .O(N__7579),
            .I(\uu2.r_addrZ0Z_7 ));
    CascadeMux I__785 (
            .O(N__7572),
            .I(N__7568));
    InMux I__784 (
            .O(N__7571),
            .I(N__7565));
    InMux I__783 (
            .O(N__7568),
            .I(N__7560));
    LocalMux I__782 (
            .O(N__7565),
            .I(N__7557));
    InMux I__781 (
            .O(N__7564),
            .I(N__7552));
    InMux I__780 (
            .O(N__7563),
            .I(N__7552));
    LocalMux I__779 (
            .O(N__7560),
            .I(\uu2.r_addrZ0Z_6 ));
    Odrv4 I__778 (
            .O(N__7557),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__777 (
            .O(N__7552),
            .I(\uu2.r_addrZ0Z_6 ));
    InMux I__776 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__775 (
            .O(N__7542),
            .I(N__7539));
    Odrv4 I__774 (
            .O(N__7539),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    InMux I__773 (
            .O(N__7536),
            .I(N__7533));
    LocalMux I__772 (
            .O(N__7533),
            .I(N__7530));
    Odrv4 I__771 (
            .O(N__7530),
            .I(vbuf_tx_data_5));
    InMux I__770 (
            .O(N__7527),
            .I(N__7524));
    LocalMux I__769 (
            .O(N__7524),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__768 (
            .O(N__7521),
            .I(N__7518));
    LocalMux I__767 (
            .O(N__7518),
            .I(N__7515));
    Odrv4 I__766 (
            .O(N__7515),
            .I(vbuf_tx_data_6));
    InMux I__765 (
            .O(N__7512),
            .I(N__7509));
    LocalMux I__764 (
            .O(N__7509),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__763 (
            .O(N__7506),
            .I(N__7503));
    LocalMux I__762 (
            .O(N__7503),
            .I(N__7500));
    Odrv4 I__761 (
            .O(N__7500),
            .I(vbuf_tx_data_7));
    InMux I__760 (
            .O(N__7497),
            .I(N__7494));
    LocalMux I__759 (
            .O(N__7494),
            .I(N__7491));
    Odrv4 I__758 (
            .O(N__7491),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__757 (
            .O(N__7488),
            .I(N__7485));
    LocalMux I__756 (
            .O(N__7485),
            .I(N__7481));
    CEMux I__755 (
            .O(N__7484),
            .I(N__7478));
    Span4Mux_v I__754 (
            .O(N__7481),
            .I(N__7475));
    LocalMux I__753 (
            .O(N__7478),
            .I(N__7472));
    Span4Mux_s1_h I__752 (
            .O(N__7475),
            .I(N__7469));
    Span4Mux_v I__751 (
            .O(N__7472),
            .I(N__7466));
    Odrv4 I__750 (
            .O(N__7469),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__749 (
            .O(N__7466),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    CEMux I__748 (
            .O(N__7461),
            .I(N__7458));
    LocalMux I__747 (
            .O(N__7458),
            .I(N__7454));
    CEMux I__746 (
            .O(N__7457),
            .I(N__7451));
    Span4Mux_v I__745 (
            .O(N__7454),
            .I(N__7448));
    LocalMux I__744 (
            .O(N__7451),
            .I(N__7445));
    Odrv4 I__743 (
            .O(N__7448),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    Odrv12 I__742 (
            .O(N__7445),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    InMux I__741 (
            .O(N__7440),
            .I(N__7437));
    LocalMux I__740 (
            .O(N__7437),
            .I(\uu2.r_data_wire_0 ));
    InMux I__739 (
            .O(N__7434),
            .I(N__7431));
    LocalMux I__738 (
            .O(N__7431),
            .I(vbuf_tx_data_0));
    InMux I__737 (
            .O(N__7428),
            .I(N__7425));
    LocalMux I__736 (
            .O(N__7425),
            .I(N__7422));
    Odrv4 I__735 (
            .O(N__7422),
            .I(\uu2.r_data_wire_1 ));
    InMux I__734 (
            .O(N__7419),
            .I(N__7416));
    LocalMux I__733 (
            .O(N__7416),
            .I(vbuf_tx_data_1));
    InMux I__732 (
            .O(N__7413),
            .I(N__7410));
    LocalMux I__731 (
            .O(N__7410),
            .I(\uu2.r_data_wire_2 ));
    InMux I__730 (
            .O(N__7407),
            .I(N__7404));
    LocalMux I__729 (
            .O(N__7404),
            .I(vbuf_tx_data_2));
    InMux I__728 (
            .O(N__7401),
            .I(N__7398));
    LocalMux I__727 (
            .O(N__7398),
            .I(\uu2.r_data_wire_3 ));
    InMux I__726 (
            .O(N__7395),
            .I(N__7392));
    LocalMux I__725 (
            .O(N__7392),
            .I(vbuf_tx_data_3));
    InMux I__724 (
            .O(N__7389),
            .I(N__7386));
    LocalMux I__723 (
            .O(N__7386),
            .I(\uu2.r_data_wire_5 ));
    InMux I__722 (
            .O(N__7383),
            .I(N__7380));
    LocalMux I__721 (
            .O(N__7380),
            .I(\uu2.r_data_wire_6 ));
    InMux I__720 (
            .O(N__7377),
            .I(N__7374));
    LocalMux I__719 (
            .O(N__7374),
            .I(\uu2.r_data_wire_7 ));
    CascadeMux I__718 (
            .O(N__7371),
            .I(N__7368));
    InMux I__717 (
            .O(N__7368),
            .I(N__7362));
    InMux I__716 (
            .O(N__7367),
            .I(N__7362));
    LocalMux I__715 (
            .O(N__7362),
            .I(N__7359));
    Odrv4 I__714 (
            .O(N__7359),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    InMux I__713 (
            .O(N__7356),
            .I(N__7351));
    InMux I__712 (
            .O(N__7355),
            .I(N__7348));
    InMux I__711 (
            .O(N__7354),
            .I(N__7345));
    LocalMux I__710 (
            .O(N__7351),
            .I(N__7339));
    LocalMux I__709 (
            .O(N__7348),
            .I(N__7339));
    LocalMux I__708 (
            .O(N__7345),
            .I(N__7336));
    InMux I__707 (
            .O(N__7344),
            .I(N__7333));
    Odrv12 I__706 (
            .O(N__7339),
            .I(\uu0.un66_ci ));
    Odrv4 I__705 (
            .O(N__7336),
            .I(\uu0.un66_ci ));
    LocalMux I__704 (
            .O(N__7333),
            .I(\uu0.un66_ci ));
    CascadeMux I__703 (
            .O(N__7326),
            .I(N__7322));
    InMux I__702 (
            .O(N__7325),
            .I(N__7319));
    InMux I__701 (
            .O(N__7322),
            .I(N__7316));
    LocalMux I__700 (
            .O(N__7319),
            .I(N__7311));
    LocalMux I__699 (
            .O(N__7316),
            .I(N__7311));
    Odrv4 I__698 (
            .O(N__7311),
            .I(\uu0.un88_ci_3 ));
    CascadeMux I__697 (
            .O(N__7308),
            .I(\uu0.un66_ci_cascade_ ));
    InMux I__696 (
            .O(N__7305),
            .I(N__7301));
    InMux I__695 (
            .O(N__7304),
            .I(N__7296));
    LocalMux I__694 (
            .O(N__7301),
            .I(N__7293));
    InMux I__693 (
            .O(N__7300),
            .I(N__7288));
    InMux I__692 (
            .O(N__7299),
            .I(N__7288));
    LocalMux I__691 (
            .O(N__7296),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv12 I__690 (
            .O(N__7293),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__689 (
            .O(N__7288),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__688 (
            .O(N__7281),
            .I(N__7276));
    InMux I__687 (
            .O(N__7280),
            .I(N__7271));
    InMux I__686 (
            .O(N__7279),
            .I(N__7271));
    LocalMux I__685 (
            .O(N__7276),
            .I(N__7268));
    LocalMux I__684 (
            .O(N__7271),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv12 I__683 (
            .O(N__7268),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__682 (
            .O(N__7263),
            .I(N__7257));
    InMux I__681 (
            .O(N__7262),
            .I(N__7247));
    InMux I__680 (
            .O(N__7261),
            .I(N__7247));
    InMux I__679 (
            .O(N__7260),
            .I(N__7247));
    InMux I__678 (
            .O(N__7257),
            .I(N__7247));
    InMux I__677 (
            .O(N__7256),
            .I(N__7244));
    LocalMux I__676 (
            .O(N__7247),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__675 (
            .O(N__7244),
            .I(\uu0.l_countZ0Z_1 ));
    InMux I__674 (
            .O(N__7239),
            .I(N__7236));
    LocalMux I__673 (
            .O(N__7236),
            .I(N__7233));
    Odrv4 I__672 (
            .O(N__7233),
            .I(\uu0.un4_l_count_12 ));
    CascadeMux I__671 (
            .O(N__7230),
            .I(N__7227));
    InMux I__670 (
            .O(N__7227),
            .I(N__7223));
    CascadeMux I__669 (
            .O(N__7226),
            .I(N__7220));
    LocalMux I__668 (
            .O(N__7223),
            .I(N__7217));
    InMux I__667 (
            .O(N__7220),
            .I(N__7214));
    Odrv4 I__666 (
            .O(N__7217),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__665 (
            .O(N__7214),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__664 (
            .O(N__7209),
            .I(\uu0.un154_ci_9_cascade_ ));
    InMux I__663 (
            .O(N__7206),
            .I(N__7196));
    InMux I__662 (
            .O(N__7205),
            .I(N__7196));
    InMux I__661 (
            .O(N__7204),
            .I(N__7196));
    InMux I__660 (
            .O(N__7203),
            .I(N__7193));
    LocalMux I__659 (
            .O(N__7196),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__658 (
            .O(N__7193),
            .I(\uu0.l_countZ0Z_14 ));
    CascadeMux I__657 (
            .O(N__7188),
            .I(N__7183));
    InMux I__656 (
            .O(N__7187),
            .I(N__7178));
    InMux I__655 (
            .O(N__7186),
            .I(N__7178));
    InMux I__654 (
            .O(N__7183),
            .I(N__7175));
    LocalMux I__653 (
            .O(N__7178),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__652 (
            .O(N__7175),
            .I(\uu0.l_countZ0Z_15 ));
    InMux I__651 (
            .O(N__7170),
            .I(N__7164));
    InMux I__650 (
            .O(N__7169),
            .I(N__7161));
    InMux I__649 (
            .O(N__7168),
            .I(N__7158));
    InMux I__648 (
            .O(N__7167),
            .I(N__7155));
    LocalMux I__647 (
            .O(N__7164),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__646 (
            .O(N__7161),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__645 (
            .O(N__7158),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__644 (
            .O(N__7155),
            .I(\uu0.l_countZ0Z_4 ));
    CascadeMux I__643 (
            .O(N__7146),
            .I(\uu0.un4_l_count_13_cascade_ ));
    CascadeMux I__642 (
            .O(N__7143),
            .I(\uu0.un4_l_count_0_cascade_ ));
    IoInMux I__641 (
            .O(N__7140),
            .I(N__7137));
    LocalMux I__640 (
            .O(N__7137),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__639 (
            .O(N__7134),
            .I(\uu0.un4_l_count_11_cascade_ ));
    InMux I__638 (
            .O(N__7131),
            .I(N__7128));
    LocalMux I__637 (
            .O(N__7128),
            .I(\uu0.un4_l_count_16 ));
    InMux I__636 (
            .O(N__7125),
            .I(N__7118));
    InMux I__635 (
            .O(N__7124),
            .I(N__7118));
    InMux I__634 (
            .O(N__7123),
            .I(N__7115));
    LocalMux I__633 (
            .O(N__7118),
            .I(N__7112));
    LocalMux I__632 (
            .O(N__7115),
            .I(\uu0.l_countZ0Z_7 ));
    Odrv4 I__631 (
            .O(N__7112),
            .I(\uu0.l_countZ0Z_7 ));
    CascadeMux I__630 (
            .O(N__7107),
            .I(\uu0.un88_ci_3_cascade_ ));
    CascadeMux I__629 (
            .O(N__7104),
            .I(N__7101));
    InMux I__628 (
            .O(N__7101),
            .I(N__7098));
    LocalMux I__627 (
            .O(N__7098),
            .I(\uu0.un99_ci_0 ));
    CascadeMux I__626 (
            .O(N__7095),
            .I(\uu0.un187_ci_1_cascade_ ));
    InMux I__625 (
            .O(N__7092),
            .I(N__7089));
    LocalMux I__624 (
            .O(N__7089),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__623 (
            .O(N__7086),
            .I(N__7083));
    LocalMux I__622 (
            .O(N__7083),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__621 (
            .O(N__7080),
            .I(N__7077));
    LocalMux I__620 (
            .O(N__7077),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__619 (
            .O(N__7074),
            .I(N__7071));
    LocalMux I__618 (
            .O(N__7071),
            .I(vbuf_tx_data_4));
    InMux I__617 (
            .O(N__7068),
            .I(N__7065));
    LocalMux I__616 (
            .O(N__7065),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__615 (
            .O(N__7062),
            .I(N__7059));
    LocalMux I__614 (
            .O(N__7059),
            .I(N__7056));
    Span4Mux_v I__613 (
            .O(N__7056),
            .I(N__7053));
    Odrv4 I__612 (
            .O(N__7053),
            .I(\uu2.r_data_wire_4 ));
    InMux I__611 (
            .O(N__7050),
            .I(N__7047));
    LocalMux I__610 (
            .O(N__7047),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__609 (
            .O(N__7044),
            .I(N__7041));
    LocalMux I__608 (
            .O(N__7041),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__607 (
            .O(N__7038),
            .I(N__7035));
    LocalMux I__606 (
            .O(N__7035),
            .I(N__7032));
    IoSpan4Mux I__605 (
            .O(N__7032),
            .I(N__7029));
    Span4Mux_s0_h I__604 (
            .O(N__7029),
            .I(N__7026));
    Odrv4 I__603 (
            .O(N__7026),
            .I(o_serial_data_c));
    IoInMux I__602 (
            .O(N__7023),
            .I(N__7020));
    LocalMux I__601 (
            .O(N__7020),
            .I(N__7017));
    IoSpan4Mux I__600 (
            .O(N__7017),
            .I(N__7014));
    Odrv4 I__599 (
            .O(N__7014),
            .I(clk_in_c));
    INV \INVuu2.bitmap_58C  (
            .O(\INVuu2.bitmap_58C_net ),
            .I(N__18484));
    INV \INVuu2.w_addr_displaying_7_rep1C  (
            .O(\INVuu2.w_addr_displaying_7_rep1C_net ),
            .I(N__18492));
    INV \INVuu2.w_addr_displaying_ness_6C  (
            .O(\INVuu2.w_addr_displaying_ness_6C_net ),
            .I(N__18499));
    INV \INVuu2.bitmap_168C  (
            .O(\INVuu2.bitmap_168C_net ),
            .I(N__18504));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__18507));
    INV \INVuu2.bitmap_180C  (
            .O(\INVuu2.bitmap_180C_net ),
            .I(N__18460));
    INV \INVuu2.bitmap_34C  (
            .O(\INVuu2.bitmap_34C_net ),
            .I(N__18467));
    INV \INVuu2.w_addr_displaying_4_rep1C  (
            .O(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .I(N__18483));
    INV \INVuu2.bitmap_75C  (
            .O(\INVuu2.bitmap_75C_net ),
            .I(N__18498));
    INV \INVuu2.bitmap_162C  (
            .O(\INVuu2.bitmap_162C_net ),
            .I(N__18503));
    INV \INVuu2.w_addr_displaying_3_rep1_nesrC  (
            .O(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .I(N__18459));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__18466));
    INV \INVuu2.w_addr_displaying_1C  (
            .O(\INVuu2.w_addr_displaying_1C_net ),
            .I(N__18475));
    INV \INVuu2.bitmap_90C  (
            .O(\INVuu2.bitmap_90C_net ),
            .I(N__18497));
    INV \INVuu2.w_addr_displaying_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .I(N__18448));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__18477));
    INV \INVuu2.w_addr_displaying_0C  (
            .O(\INVuu2.w_addr_displaying_0C_net ),
            .I(N__18474));
    INV \INVuu2.w_addr_user_nesr_0C  (
            .O(\INVuu2.w_addr_user_nesr_0C_net ),
            .I(N__18482));
    INV \INVuu2.w_addr_user_1C  (
            .O(\INVuu2.w_addr_user_1C_net ),
            .I(N__18473));
    INV \INVuu2.w_addr_user_8C  (
            .O(\INVuu2.w_addr_user_8C_net ),
            .I(N__18489));
    INV \INVuu2.bitmap_111C  (
            .O(\INVuu2.bitmap_111C_net ),
            .I(N__18472));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__18501));
    INV \INVuu2.r_data_reg_4C  (
            .O(\INVuu2.r_data_reg_4C_net ),
            .I(N__18505));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__10533),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__7140),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__10362),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_1_5_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7062),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_4C_net ),
            .ce(N__7461),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_1_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_1_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_1_6_0  (
            .in0(N__8883),
            .in1(N__7092),
            .in2(_gnd_net_),
            .in3(N__7434),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.shifter_0_LC_1_6_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_1_6_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__7050),
            .in2(_gnd_net_),
            .in3(N__8881),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.uart_tx_LC_1_6_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_1_6_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_1_6_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_1_6_2  (
            .in0(N__8882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7044),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.shifter_2_LC_1_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_1_6_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_1_6_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_1_6_3  (
            .in0(N__7086),
            .in1(N__8884),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.shifter_3_LC_1_6_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_1_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_1_6_4  (
            .in0(N__8885),
            .in1(N__7080),
            .in2(_gnd_net_),
            .in3(N__7407),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.shifter_4_LC_1_6_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_1_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_1_6_5  (
            .in0(N__7068),
            .in1(N__8886),
            .in2(_gnd_net_),
            .in3(N__7395),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \buart.Z_tx.shifter_5_LC_1_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_1_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_1_6_6  (
            .in0(N__8887),
            .in1(N__7527),
            .in2(_gnd_net_),
            .in3(N__7074),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18500),
            .ce(N__7484),
            .sr(N__18700));
    defparam \uu0.l_count_13_LC_1_7_1 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_7_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_7_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_13_LC_1_7_1  (
            .in0(N__7895),
            .in1(N__9721),
            .in2(N__7767),
            .in3(N__7824),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18493),
            .ce(N__8195),
            .sr(N__18698));
    defparam \uu0.l_count_7_LC_1_7_2 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_1_7_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_1_7_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_7_LC_1_7_2  (
            .in0(N__9722),
            .in1(N__7356),
            .in2(N__7104),
            .in3(N__7123),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18493),
            .ce(N__8195),
            .sr(N__18698));
    defparam \uu0.l_count_12_LC_1_7_6 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_7_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_12_LC_1_7_6  (
            .in0(N__9720),
            .in1(N__7896),
            .in2(N__7797),
            .in3(N__7812),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18493),
            .ce(N__8195),
            .sr(N__18698));
    defparam \uu0.l_count_16_LC_1_8_2 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_1_8_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_16_LC_1_8_2  (
            .in0(N__7897),
            .in1(N__9719),
            .in2(N__7845),
            .in3(N__8067),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18487),
            .ce(N__8193),
            .sr(N__18697));
    defparam \uu0.l_count_8_LC_1_8_3 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_8_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_count_8_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__7898),
            .in2(_gnd_net_),
            .in3(N__8754),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18487),
            .ce(N__8193),
            .sr(N__18697));
    defparam \uu0.l_count_5_LC_1_8_4 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_1_8_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu0.l_count_5_LC_1_8_4  (
            .in0(N__7280),
            .in1(N__7355),
            .in2(_gnd_net_),
            .in3(N__7170),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18487),
            .ce(N__8193),
            .sr(N__18697));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__7168),
            .in2(_gnd_net_),
            .in3(N__7279),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(\uu0.un88_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_8_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_8_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7107),
            .in3(N__7305),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_1_8_7 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_1_8_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_1_8_7  (
            .in0(N__7988),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7977),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_10_LC_1_9_1 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_9_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu0.l_count_10_LC_1_9_1  (
            .in0(N__8750),
            .in1(N__7894),
            .in2(N__8786),
            .in3(N__8710),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18479),
            .ce(N__8192),
            .sr(N__18699));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_9_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_9_2  (
            .in0(N__7205),
            .in1(N__7788),
            .in2(_gnd_net_),
            .in3(N__8042),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_9_3 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_9_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_15_LC_1_9_3  (
            .in0(N__7890),
            .in1(N__9704),
            .in2(N__7095),
            .in3(N__7187),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18479),
            .ce(N__8192),
            .sr(N__18699));
    defparam \uu0.l_count_14_LC_1_9_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_9_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_14_LC_1_9_4  (
            .in0(N__7206),
            .in1(N__8043),
            .in2(N__7899),
            .in3(N__7789),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18479),
            .ce(N__8192),
            .sr(N__18699));
    defparam \uu0.l_count_4_LC_1_9_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_9_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \uu0.l_count_4_LC_1_9_5  (
            .in0(N__7354),
            .in1(N__9705),
            .in2(_gnd_net_),
            .in3(N__7169),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18479),
            .ce(N__8192),
            .sr(N__18699));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_9_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_9_6  (
            .in0(N__8709),
            .in1(N__8779),
            .in2(N__7922),
            .in3(N__8749),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_9_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_9_7  (
            .in0(N__8041),
            .in1(N__7186),
            .in2(N__7209),
            .in3(N__7204),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIGTCU_15_LC_1_10_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_10_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu0.l_count_RNIGTCU_15_LC_1_10_0  (
            .in0(N__8778),
            .in1(N__7203),
            .in2(N__7188),
            .in3(N__7167),
            .lcout(),
            .ltout(\uu0.un4_l_count_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_10_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_15_LC_1_10_1  (
            .in0(N__7239),
            .in1(N__7131),
            .in2(N__7146),
            .in3(N__8019),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_2 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_2 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__9996),
            .in2(N__7143),
            .in3(N__10007),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_1_10_3 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_1_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.sec_clkD_LC_1_10_3  (
            .in0(N__9663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.sec_clkDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18471),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_10_4 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_10_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_1_10_4  (
            .in0(N__8708),
            .in1(N__7124),
            .in2(N__8229),
            .in3(N__7939),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNIOIDD2_18_LC_1_10_5  (
            .in0(N__7915),
            .in1(N__8207),
            .in2(N__7134),
            .in3(N__7299),
            .lcout(\uu0.un4_l_count_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_10_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_10_7  (
            .in0(N__7125),
            .in1(N__7344),
            .in2(N__7326),
            .in3(N__7300),
            .lcout(\uu0.un110_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_11_1 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_11_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_2_LC_1_11_1  (
            .in0(N__8097),
            .in1(N__7262),
            .in2(_gnd_net_),
            .in3(N__8133),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18462),
            .ce(N__8194),
            .sr(N__18701));
    defparam \uu0.l_count_1_LC_1_11_2 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_11_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_11_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_1_11_2  (
            .in0(N__7261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8096),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18462),
            .ce(N__8194),
            .sr(N__18701));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_3  (
            .in0(N__8094),
            .in1(N__7260),
            .in2(_gnd_net_),
            .in3(N__8132),
            .lcout(\uu0.un55_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_0_LC_1_11_4 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_11_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_11_4  (
            .in0(N__9699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8095),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18462),
            .ce(N__8194),
            .sr(N__18701));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_6  (
            .in0(N__8131),
            .in1(N__7940),
            .in2(N__7263),
            .in3(N__8093),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_6_LC_1_11_7 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_1_11_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_6_LC_1_11_7  (
            .in0(N__7325),
            .in1(N__9700),
            .in2(N__7308),
            .in3(N__7304),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18462),
            .ce(N__8194),
            .sr(N__18701));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_1_12_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_1_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__8869),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_12_6 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_12_6  (
            .in0(N__8150),
            .in1(N__7281),
            .in2(N__8175),
            .in3(N__7256),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_2_4_0 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_2_4_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_8_LC_2_4_0  (
            .in0(N__7545),
            .in1(N__7367),
            .in2(N__7226),
            .in3(N__7714),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18506),
            .ce(N__7659),
            .sr(N__18689));
    defparam \uu2.r_addr_esr_3_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_2_4_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_2_4_4  (
            .in0(N__15893),
            .in1(N__15768),
            .in2(N__7630),
            .in3(N__15835),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18506),
            .ce(N__7659),
            .sr(N__18689));
    defparam \uu2.r_addr_esr_7_LC_2_4_7 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_2_4_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_2_4_7  (
            .in0(N__7715),
            .in1(N__7591),
            .in2(N__7371),
            .in3(N__7571),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18506),
            .ce(N__7659),
            .sr(N__18689));
    defparam \uu2.r_data_reg_0_LC_2_5_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_0_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7440),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_5_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_1_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7428),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_2_LC_2_5_2  (
            .in0(N__7413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_5_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_3_LC_2_5_3  (
            .in0(N__7401),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_5_LC_2_5_5  (
            .in0(N__7389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7383),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_5_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7377),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7457),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__7741),
            .in2(_gnd_net_),
            .in3(N__7684),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_6_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_6_4  (
            .in0(N__15889),
            .in1(N__15754),
            .in2(N__7634),
            .in3(N__15834),
            .lcout(\uu2.un404_ci ),
            .ltout(\uu2.un404_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_2_6_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_2_6_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_6_LC_2_6_5  (
            .in0(N__7564),
            .in1(N__7742),
            .in2(N__7602),
            .in3(N__7685),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18494),
            .ce(N__7655),
            .sr(N__18688));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_6_6 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__7595),
            .in2(_gnd_net_),
            .in3(N__7563),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI83ID7_8_LC_2_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI83ID7_8_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI83ID7_8_LC_2_6_7 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI83ID7_8_LC_2_6_7  (
            .in0(N__9152),
            .in1(N__14682),
            .in2(N__12810),
            .in3(N__11844),
            .lcout(\uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_6_LC_2_7_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_7_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_7_0  (
            .in0(N__7512),
            .in1(N__8872),
            .in2(_gnd_net_),
            .in3(N__7536),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18488),
            .ce(N__7488),
            .sr(N__18742));
    defparam \buart.Z_tx.shifter_7_LC_2_7_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_7_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_7_1  (
            .in0(N__8873),
            .in1(N__7497),
            .in2(_gnd_net_),
            .in3(N__7521),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18488),
            .ce(N__7488),
            .sr(N__18742));
    defparam \buart.Z_tx.shifter_8_LC_2_7_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_7_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_7_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__8871),
            .in2(_gnd_net_),
            .in3(N__7506),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18488),
            .ce(N__7488),
            .sr(N__18742));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_7_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_7_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_2_7_3  (
            .in0(N__7956),
            .in1(N__7971),
            .in2(_gnd_net_),
            .in3(N__18741),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIMBBL2_7_LC_2_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIMBBL2_7_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIMBBL2_7_LC_2_7_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIMBBL2_7_LC_2_7_4  (
            .in0(N__15398),
            .in1(N__15197),
            .in2(_gnd_net_),
            .in3(N__15339),
            .lcout(\uu2.N_15_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__7823),
            .in2(_gnd_net_),
            .in3(N__7810),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_6  (
            .in0(N__7811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7793),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_2_7_7 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_7_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__7758),
            .in2(_gnd_net_),
            .in3(N__9659),
            .lcout(oneSecStrb_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_5_LC_2_8_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_2_8_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_5_LC_2_8_0  (
            .in0(N__15788),
            .in1(N__7683),
            .in2(N__7716),
            .in3(N__7737),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \uu2.r_addr_4_LC_2_8_1 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_2_8_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_2_8_1  (
            .in0(N__7682),
            .in1(N__7710),
            .in2(_gnd_net_),
            .in3(N__15787),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_8_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_8_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_2_8_2  (
            .in0(N__15785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18747),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_0_LC_2_8_3 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_2_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.r_addr_0_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__15824),
            .in2(_gnd_net_),
            .in3(N__15786),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_2_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_2_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_1_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__9599),
            .in2(_gnd_net_),
            .in3(N__9578),
            .lcout(\Lab_UT.alarmchar10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_2_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_2_8_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_2_8_5 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_2_LC_2_8_5  (
            .in0(N__9579),
            .in1(_gnd_net_),
            .in2(N__9603),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmchar10_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \uu2.trig_rd_det_0_LC_2_8_6 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_2_8_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__10074),
            .in2(_gnd_net_),
            .in3(N__8670),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \uu2.trig_rd_det_1_LC_2_8_7 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_2_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7989),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18480),
            .ce(),
            .sr(N__18687));
    defparam \uu2.bitmap_111_LC_2_9_0 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_2_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9652),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__18648));
    defparam \uu2.vram_rd_clk_det_0_LC_2_9_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_2_9_1 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10069),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__18648));
    defparam \uu2.vram_rd_clk_det_1_LC_2_9_2 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_2_9_2 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7970),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__18648));
    defparam \uu0.l_count_3_LC_2_10_1 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_2_10_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \uu0.l_count_3_LC_2_10_1  (
            .in0(N__7947),
            .in1(N__9703),
            .in2(_gnd_net_),
            .in3(N__7941),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18463),
            .ce(N__8196),
            .sr(N__18702));
    defparam \uu0.l_count_9_LC_2_10_2 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_2_10_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_9_LC_2_10_2  (
            .in0(N__7887),
            .in1(N__8756),
            .in2(_gnd_net_),
            .in3(N__8714),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18463),
            .ce(N__8196),
            .sr(N__18702));
    defparam \uu0.l_count_17_LC_2_10_3 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_10_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_10_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_17_LC_2_10_3  (
            .in0(N__8228),
            .in1(N__7840),
            .in2(N__8073),
            .in3(N__7889),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18463),
            .ce(N__8196),
            .sr(N__18702));
    defparam \uu0.l_count_11_LC_2_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_2_10_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_2_10_5 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uu0.l_count_11_LC_2_10_5  (
            .in0(N__8685),
            .in1(N__9701),
            .in2(N__7923),
            .in3(N__7888),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18463),
            .ce(N__8196),
            .sr(N__18702));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_10_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_10_6  (
            .in0(N__7886),
            .in1(N__8069),
            .in2(N__7844),
            .in3(N__8227),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_10_7 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_10_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_10_7 .LUT_INIT=16'b0001001000010010;
    LogicCell40 \uu0.l_count_18_LC_2_10_7  (
            .in0(N__8208),
            .in1(N__9702),
            .in2(N__8211),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18463),
            .ce(N__8196),
            .sr(N__18702));
    defparam \uu0.delay_line_0_LC_2_11_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_2_11_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_2_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_2_11_0  (
            .in0(N__8173),
            .in1(N__8151),
            .in2(N__8013),
            .in3(N__8112),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18456),
            .ce(),
            .sr(N__18703));
    defparam \uu0.l_precount_3_LC_2_11_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_2_11_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_2_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_precount_3_LC_2_11_1  (
            .in0(N__8114),
            .in1(N__8012),
            .in2(N__8157),
            .in3(N__8174),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18456),
            .ce(),
            .sr(N__18703));
    defparam \uu0.l_precount_1_LC_2_11_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_2_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_2_11_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_precount_1_LC_2_11_3  (
            .in0(N__8152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8010),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18456),
            .ce(),
            .sr(N__18703));
    defparam \uu0.l_precount_2_LC_2_11_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_2_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_2_11_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_2_11_4  (
            .in0(N__8011),
            .in1(N__8153),
            .in2(_gnd_net_),
            .in3(N__8113),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18456),
            .ce(),
            .sr(N__18703));
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_2_11_5 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_2_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI3Q7K1_2_LC_2_11_5  (
            .in0(N__8755),
            .in1(N__8130),
            .in2(N__8115),
            .in3(N__8092),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNIO2782_16_LC_2_11_6  (
            .in0(N__8005),
            .in1(N__8068),
            .in2(N__8046),
            .in3(N__8040),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_0_LC_2_11_7 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_2_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8009),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18456),
            .ce(),
            .sr(N__18703));
    defparam \buart.Z_tx.bitcount_0_LC_2_12_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_2_12_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_2_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_2_12_0  (
            .in0(N__8870),
            .in1(N__8288),
            .in2(_gnd_net_),
            .in3(N__8328),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18449),
            .ce(),
            .sr(N__18704));
    defparam \buart.Z_tx.bitcount_1_LC_2_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_2_13_0 .LUT_INIT=16'b1111110011110110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_2_13_0  (
            .in0(N__8325),
            .in1(N__8304),
            .in2(N__8888),
            .in3(N__8287),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18442),
            .ce(),
            .sr(N__18706));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_13_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_13_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_2_13_1  (
            .in0(N__8303),
            .in1(N__8256),
            .in2(N__8289),
            .in3(N__8324),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_2_13_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_2_13_2 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_2_13_2  (
            .in0(N__8326),
            .in1(N__8889),
            .in2(N__8346),
            .in3(N__8343),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18442),
            .ce(),
            .sr(N__18706));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_13_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__8282),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_13_4 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_13_4  (
            .in0(N__8254),
            .in1(N__8301),
            .in2(N__8331),
            .in3(N__9024),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_13_5 .LUT_INIT=16'b1110111100010000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_2_13_5  (
            .in0(N__8302),
            .in1(N__8283),
            .in2(N__8262),
            .in3(N__8255),
            .lcout(),
            .ltout(\buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_2_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_2_13_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_2_13_6  (
            .in0(N__8874),
            .in1(_gnd_net_),
            .in2(N__8259),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18442),
            .ce(),
            .sr(N__18706));
    defparam \Lab_UT.alarmchar_5_LC_4_3_2 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_5_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_5_LC_4_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.alarmchar_5_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8244),
            .lcout(\Lab_UT.alarmcharZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18502),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNO_0_8_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNO_0_8_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNO_0_8_LC_4_4_1 .LUT_INIT=16'b0110001100110011;
    LogicCell40 \uu2.w_addr_user_RNO_0_8_LC_4_4_1  (
            .in0(N__9391),
            .in1(N__8368),
            .in2(N__10255),
            .in3(N__9376),
            .lcout(\uu2.N_61_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_4_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_4_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_4_4_7  (
            .in0(N__14529),
            .in1(N__12372),
            .in2(N__9329),
            .in3(N__14396),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_5_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_4_5_0  (
            .in0(N__14527),
            .in1(N__15198),
            .in2(N__9378),
            .in3(N__14395),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_1  (
            .in0(N__14394),
            .in1(N__14528),
            .in2(N__8370),
            .in3(N__14668),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIK9E4_2_LC_4_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIK9E4_2_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIK9E4_2_LC_4_5_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIK9E4_2_LC_4_5_3  (
            .in0(N__12148),
            .in1(N__10306),
            .in2(_gnd_net_),
            .in3(N__10147),
            .lcout(\uu2.N_102 ),
            .ltout(\uu2.N_102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIQ6EA_5_LC_4_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIQ6EA_5_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIQ6EA_5_LC_4_5_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.w_addr_user_RNIQ6EA_5_LC_4_5_4  (
            .in0(N__9233),
            .in1(N__8513),
            .in2(N__8382),
            .in3(N__9324),
            .lcout(\uu2.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_8_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_8_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_8_LC_4_5_5 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \uu2.w_addr_user_8_LC_4_5_5  (
            .in0(N__8367),
            .in1(N__9285),
            .in2(N__8379),
            .in3(N__8550),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_8C_net ),
            .ce(),
            .sr(N__18652));
    defparam \uu2.w_addr_user_RNO_0_5_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNO_0_5_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNO_0_5_LC_4_5_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \uu2.w_addr_user_RNO_0_5_LC_4_5_6  (
            .in0(N__9346),
            .in1(N__9234),
            .in2(_gnd_net_),
            .in3(N__9325),
            .lcout(\uu2.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI86V6_2_LC_4_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI86V6_2_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI86V6_2_LC_4_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI86V6_2_LC_4_5_7  (
            .in0(N__8512),
            .in1(N__9372),
            .in2(N__8369),
            .in3(N__10146),
            .lcout(\uu2.w_addr_user_3_i_a2_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIR7FF7_6_LC_4_6_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIR7FF7_6_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIR7FF7_6_LC_4_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_user_nesr_RNIR7FF7_6_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__10357),
            .in2(_gnd_net_),
            .in3(N__8544),
            .lcout(\uu2.un28_w_addr_user_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_6_LC_4_6_1 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_6_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_6_LC_4_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.alarmchar_6_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8487),
            .lcout(\Lab_UT.alarmcharZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18481),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_6_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_6_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_4_6_2  (
            .in0(N__14375),
            .in1(N__14504),
            .in2(N__8517),
            .in3(N__15578),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI2UTD_1_LC_4_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI2UTD_1_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI2UTD_1_LC_4_6_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.w_addr_user_RNI2UTD_1_LC_4_6_3  (
            .in0(N__8469),
            .in1(N__12142),
            .in2(N__10305),
            .in3(N__8418),
            .lcout(\uu2.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_4  (
            .in0(N__13944),
            .in1(N__11085),
            .in2(N__8448),
            .in3(N__10950),
            .lcout(),
            .ltout(\uu2.mem0.g1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_6_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_6_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_6_5  (
            .in0(N__10485),
            .in1(N__8454),
            .in2(N__8463),
            .in3(N__9432),
            .lcout(\uu2.mem0.N_63_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_6 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_6  (
            .in0(N__11073),
            .in1(N__13959),
            .in2(N__8447),
            .in3(N__9528),
            .lcout(\uu2.mem0.G_17_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_4_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_4_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dispString.rdy_RNIGIDK3_LC_4_6_7  (
            .in0(N__14503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14374),
            .lcout(N_72_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_4_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_4_7_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_4_7_1  (
            .in0(N__14462),
            .in1(N__12474),
            .in2(N__9240),
            .in3(N__14353),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI0FF3_4_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI0FF3_4_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI0FF3_4_LC_4_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.w_addr_user_nesr_RNI0FF3_4_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__9236),
            .in2(_gnd_net_),
            .in3(N__9308),
            .lcout(\uu2.w_addr_user_3_i_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNINEKD7_6_LC_4_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNINEKD7_6_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNINEKD7_6_LC_4_7_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \uu2.w_addr_user_nesr_RNINEKD7_6_LC_4_7_4  (
            .in0(N__9404),
            .in1(N__9259),
            .in2(N__10260),
            .in3(N__14461),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(\uu2.un28_w_addr_user_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_1_LC_4_7_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_4_7_5 .LUT_INIT=16'b0001110001001100;
    LogicCell40 \uu2.w_addr_user_1_LC_4_7_5  (
            .in0(N__9260),
            .in1(N__10301),
            .in2(N__8553),
            .in3(N__12149),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__18649));
    defparam \uu2.w_addr_user_3_LC_4_7_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_3_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_3_LC_4_7_6 .LUT_INIT=16'b0010000110101010;
    LogicCell40 \uu2.w_addr_user_3_LC_4_7_6  (
            .in0(N__9320),
            .in1(N__9261),
            .in2(N__9354),
            .in3(N__8545),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__18649));
    defparam \uu2.w_addr_user_5_LC_4_7_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_4_7_7 .LUT_INIT=16'b0101110100000010;
    LogicCell40 \uu2.w_addr_user_5_LC_4_7_7  (
            .in0(N__8546),
            .in1(N__8526),
            .in2(N__9279),
            .in3(N__8511),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__18649));
    defparam \uu2.un28_w_addr_user_i_0_a2_0_LC_4_8_0 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_LC_4_8_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a2_0_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__9524),
            .in2(_gnd_net_),
            .in3(N__9482),
            .lcout(),
            .ltout(\uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_o4_LC_4_8_1 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_o4_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_o4_LC_4_8_1 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \uu2.un28_w_addr_user_i_0_o4_LC_4_8_1  (
            .in0(N__9534),
            .in1(N__9502),
            .in2(N__8490),
            .in3(N__14328),
            .lcout(\uu2.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_2 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_4_8_2  (
            .in0(N__10659),
            .in1(N__16723),
            .in2(N__8637),
            .in3(N__16833),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18464),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_4_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_4_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__10809),
            .in2(_gnd_net_),
            .in3(N__10776),
            .lcout(\Lab_UT.alarmchar_2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_4_8_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__8624),
            .in2(_gnd_net_),
            .in3(N__8587),
            .lcout(),
            .ltout(\resetGen.reset_count_2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_4_8_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_4_8_5 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \resetGen.reset_count_4_LC_4_8_5  (
            .in0(N__10387),
            .in1(N__8598),
            .in2(N__8649),
            .in3(N__11271),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18464),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_4_LC_4_8_6 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_4_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_4_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.alarmchar_4_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8646),
            .lcout(\Lab_UT.alarmcharZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18464),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_4_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_4_8_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_3_LC_4_8_7  (
            .in0(N__9590),
            .in1(N__9569),
            .in2(_gnd_net_),
            .in3(N__10358),
            .lcout(\Lab_UT.dictrl.un1_next_alarmstate21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18464),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_4_9_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_4_9_0 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_4_9_0  (
            .in0(N__11265),
            .in1(N__10391),
            .in2(N__8571),
            .in3(N__8613),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18457),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_4_9_1 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_4_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_4_9_1  (
            .in0(N__8612),
            .in1(N__8566),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_4_9_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_4_9_2 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_3_LC_4_9_2  (
            .in0(N__11267),
            .in1(N__10390),
            .in2(N__8628),
            .in3(N__8625),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18457),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_4_9_3 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_4_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__8611),
            .in2(_gnd_net_),
            .in3(N__8565),
            .lcout(\resetGen.un241_ci ),
            .ltout(\resetGen.un241_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_4_9_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_4_9_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_4_9_4 .LUT_INIT=16'b0100010000010100;
    LogicCell40 \resetGen.reset_count_2_LC_4_9_4  (
            .in0(N__11266),
            .in1(N__8589),
            .in2(N__8592),
            .in3(N__10389),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18457),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_4_9_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_4_9_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_4_9_5 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_4_9_5  (
            .in0(N__10388),
            .in1(N__8567),
            .in2(_gnd_net_),
            .in3(N__11264),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18457),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_4_9_6 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_4_9_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_4_9_6  (
            .in0(N__10073),
            .in1(N__8669),
            .in2(N__8868),
            .in3(N__18748),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18457),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_7  (
            .in0(N__8787),
            .in1(N__8760),
            .in2(_gnd_net_),
            .in3(N__8718),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_1_LC_4_10_1 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_4_10_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_4_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_1_LC_4_10_1  (
            .in0(N__8920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8947),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18450),
            .ce(),
            .sr(N__18705));
    defparam \uu2.l_count_0_LC_4_10_2 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_4_10_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_4_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8919),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18450),
            .ce(),
            .sr(N__18705));
    defparam \uu2.l_count_7_LC_4_10_5 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_4_10_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_4_10_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.l_count_7_LC_4_10_5  (
            .in0(N__9780),
            .in1(N__10694),
            .in2(N__8979),
            .in3(N__9749),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18450),
            .ce(),
            .sr(N__18705));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_10_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_10_6  (
            .in0(N__9748),
            .in1(N__8974),
            .in2(N__10695),
            .in3(N__9779),
            .lcout(\uu2.un350_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_11_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_11_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_4_11_1  (
            .in0(N__9746),
            .in1(N__10715),
            .in2(N__8998),
            .in3(N__8912),
            .lcout(),
            .ltout(\uu2.un1_l_count_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_11_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_4_11_2  (
            .in0(N__9965),
            .in1(N__8945),
            .in2(N__8673),
            .in3(N__8958),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_11_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_4_11_3  (
            .in0(N__9747),
            .in1(N__10716),
            .in2(N__8999),
            .in3(N__8913),
            .lcout(),
            .ltout(\uu2.un1_l_count_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_4_11_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_4_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_4_11_4  (
            .in0(N__9966),
            .in1(N__8946),
            .in2(N__8652),
            .in3(N__8957),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_4_11_5 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_4_11_5 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_4_11_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uu2.l_count_4_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__10717),
            .in2(N__9003),
            .in3(N__9778),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18443),
            .ce(),
            .sr(N__18707));
    defparam \uu2.l_count_9_LC_4_11_7 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_4_11_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_4_11_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu2.l_count_9_LC_4_11_7  (
            .in0(N__9908),
            .in1(N__9923),
            .in2(N__9000),
            .in3(N__10041),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18443),
            .ce(),
            .sr(N__18707));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_4_12_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_4_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9065),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18436),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_12_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__8949),
            .in2(_gnd_net_),
            .in3(N__8922),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_12_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_4_12_2  (
            .in0(N__10738),
            .in1(N__8978),
            .in2(N__9909),
            .in3(N__10024),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_4_12_3 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_4_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_4_12_3  (
            .in0(N__9066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9041),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18436),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_12_7 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_12_7  (
            .in0(N__10025),
            .in1(N__8948),
            .in2(N__9969),
            .in3(N__8921),
            .lcout(\uu2.un306_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_4_13_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__9064),
            .in2(N__9042),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_4_13_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_4_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9087),
            .in3(N__8892),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__18431),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_4_13_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_4_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_4_13_2  (
            .in0(N__9022),
            .in1(N__9075),
            .in2(_gnd_net_),
            .in3(N__9138),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__18431),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_4_13_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_4_13_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9114),
            .in3(N__9135),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__18431),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_4_13_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_4_13_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_4_13_4  (
            .in0(N__9023),
            .in1(_gnd_net_),
            .in2(N__9126),
            .in3(N__9132),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__18431),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_4_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_4_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_4_13_5  (
            .in0(N__9101),
            .in1(N__9021),
            .in2(_gnd_net_),
            .in3(N__9129),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18431),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_4_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_4_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_4_13_6  (
            .in0(N__9122),
            .in1(N__9110),
            .in2(N__9102),
            .in3(N__9083),
            .lcout(),
            .ltout(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_4_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_4_13_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_4_13_7  (
            .in0(N__9074),
            .in1(N__9063),
            .in2(N__9045),
            .in3(N__9037),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_1_LC_5_4_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_5_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__9809),
            .in2(_gnd_net_),
            .in3(N__16685),
            .lcout(\Lab_UT.cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18490),
            .ce(),
            .sr(N__18693));
    defparam \uu2.w_addr_user_nesr_0_LC_5_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_0_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_0_LC_5_5_0 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \uu2.w_addr_user_nesr_0_LC_5_5_0  (
            .in0(N__12147),
            .in1(N__10249),
            .in2(N__9416),
            .in3(N__9280),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_0C_net ),
            .ce(N__9207),
            .sr(N__18655));
    defparam \uu2.w_addr_user_nesr_2_LC_5_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_2_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_2_LC_5_5_1 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu2.w_addr_user_nesr_2_LC_5_5_1  (
            .in0(N__9281),
            .in1(N__12146),
            .in2(N__10311),
            .in3(N__10149),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_0C_net ),
            .ce(N__9207),
            .sr(N__18655));
    defparam \uu2.w_addr_user_nesr_6_LC_5_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_6_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_6_LC_5_5_2 .LUT_INIT=16'b0000000000001001;
    LogicCell40 \uu2.w_addr_user_nesr_6_LC_5_5_2  (
            .in0(N__9392),
            .in1(N__10250),
            .in2(N__9417),
            .in3(N__9283),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_0C_net ),
            .ce(N__9207),
            .sr(N__18655));
    defparam \uu2.w_addr_user_nesr_7_LC_5_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_5_5_3 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_5_5_3  (
            .in0(N__9284),
            .in1(N__9393),
            .in2(N__10256),
            .in3(N__9377),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_0C_net ),
            .ce(N__9207),
            .sr(N__18655));
    defparam \uu2.w_addr_user_nesr_4_LC_5_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_4_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_4_LC_5_5_4 .LUT_INIT=16'b0000000010011010;
    LogicCell40 \uu2.w_addr_user_nesr_4_LC_5_5_4  (
            .in0(N__9235),
            .in1(N__9347),
            .in2(N__9330),
            .in3(N__9282),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_0C_net ),
            .ce(N__9207),
            .sr(N__18655));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_5_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_5_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_5_6_0  (
            .in0(N__9180),
            .in1(N__9507),
            .in2(_gnd_net_),
            .in3(N__11835),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIARVM2_0_LC_5_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIARVM2_0_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIARVM2_0_LC_5_6_1 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \uu2.w_addr_displaying_RNIARVM2_0_LC_5_6_1  (
            .in0(N__15639),
            .in1(N__12261),
            .in2(_gnd_net_),
            .in3(N__15717),
            .lcout(),
            .ltout(\uu2.N_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIBTS94_8_LC_5_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIBTS94_8_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIBTS94_8_LC_5_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIBTS94_8_LC_5_6_2  (
            .in0(N__14684),
            .in1(N__12075),
            .in2(N__9183),
            .in3(N__15191),
            .lcout(\uu2.N_132_mux ),
            .ltout(\uu2.N_132_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_5_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_5_6_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_5_6_3  (
            .in0(N__11836),
            .in1(_gnd_net_),
            .in2(N__9174),
            .in3(N__9483),
            .lcout(\uu2.mem0.N_94_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIREPN6_8_LC_5_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIREPN6_8_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIREPN6_8_LC_5_6_4 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIREPN6_8_LC_5_6_4  (
            .in0(N__14685),
            .in1(_gnd_net_),
            .in2(N__9159),
            .in3(N__11834),
            .lcout(\uu2.un21_w_addr_displaying_i ),
            .ltout(\uu2.un21_w_addr_displaying_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_5_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_5_6_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_0_LC_5_6_5  (
            .in0(N__15640),
            .in1(_gnd_net_),
            .in2(N__9459),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__18653));
    defparam \uu2.w_addr_displaying_fast_1_LC_5_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_1_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_1_LC_5_6_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_displaying_fast_1_LC_5_6_6  (
            .in0(N__15430),
            .in1(N__15641),
            .in2(_gnd_net_),
            .in3(N__10431),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__18653));
    defparam \uu2.w_addr_displaying_0_rep1_LC_5_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_5_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__11943),
            .in2(_gnd_net_),
            .in3(N__15429),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__18653));
    defparam \Lab_UT.bcd2segment1.m68_bm_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m68_bm_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m68_bm_LC_5_7_0 .LUT_INIT=16'b0000011100110111;
    LogicCell40 \Lab_UT.bcd2segment1.m68_bm_LC_5_7_0  (
            .in0(N__10458),
            .in1(N__16825),
            .in2(N__16722),
            .in3(N__19443),
            .lcout(\Lab_UT.bcd2segment1.m68_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_1 .LUT_INIT=16'b0010001011000100;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_5_7_1  (
            .in0(N__16826),
            .in1(N__10662),
            .in2(N__9456),
            .in3(N__16706),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18465),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_5_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_5_7_2 .LUT_INIT=16'b0101111111110011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_30_LC_5_7_2  (
            .in0(N__11176),
            .in1(N__12472),
            .in2(N__12771),
            .in3(N__12324),
            .lcout(\uu2.mem0.N_13_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_5_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_5_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIDKOL_1_LC_5_7_3  (
            .in0(N__15643),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11178),
            .lcout(\uu2.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_7_4 .LUT_INIT=16'b1111100101100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_32_LC_5_7_4  (
            .in0(N__11177),
            .in1(N__15642),
            .in2(N__10191),
            .in3(N__11976),
            .lcout(),
            .ltout(\uu2.mem0.i14_mux_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_5_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_5_7_5 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_18_LC_5_7_5  (
            .in0(N__12558),
            .in1(N__9441),
            .in2(N__9435),
            .in3(N__12618),
            .lcout(\uu2.mem0.N_8_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_5_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_5_7_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_5_7_6  (
            .in0(N__16705),
            .in1(N__16827),
            .in2(N__9426),
            .in3(N__10658),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18465),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_5_7_7  (
            .in0(N__10657),
            .in1(N__9627),
            .in2(_gnd_net_),
            .in3(N__9549),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18465),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_5_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_5_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dispString.rdy_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9810),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18458),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_5_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_5_8_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_5_8_1  (
            .in0(N__10660),
            .in1(N__9540),
            .in2(_gnd_net_),
            .in3(N__10401),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18458),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_a2_4_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a2_4_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a2_4_LC_5_8_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a2_4_LC_5_8_2  (
            .in0(N__14414),
            .in1(N__11861),
            .in2(N__10109),
            .in3(N__11041),
            .lcout(\uu2.un28_w_addr_user_i_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_5_8_3  (
            .in0(N__10661),
            .in1(N__10596),
            .in2(_gnd_net_),
            .in3(N__9618),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18458),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_8_4 .LUT_INIT=16'b0001001001001001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_47_LC_5_8_4  (
            .in0(N__12473),
            .in1(N__11164),
            .in2(N__12754),
            .in3(N__12328),
            .lcout(\uu2.mem0.g0_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_data_i_o2_4_0_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.w_data_i_o2_4_0_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_data_i_o2_4_0_LC_5_8_5 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \uu2.w_data_i_o2_4_0_LC_5_8_5  (
            .in0(N__9523),
            .in1(N__14413),
            .in2(N__9506),
            .in3(N__9481),
            .lcout(),
            .ltout(\uu2.w_data_i_o2_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_data_i_o2_0_LC_5_8_6 .C_ON=1'b0;
    defparam \uu2.w_data_i_o2_0_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_data_i_o2_0_LC_5_8_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \uu2.w_data_i_o2_0_LC_5_8_6  (
            .in0(N__10105),
            .in1(N__11860),
            .in2(N__9465),
            .in3(N__11042),
            .lcout(N_96),
            .ltout(N_96_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_data_i_0_tz_0_LC_5_8_7 .C_ON=1'b0;
    defparam \uu2.w_data_i_0_tz_0_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_data_i_0_tz_0_LC_5_8_7 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \uu2.w_data_i_0_tz_0_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9462),
            .in3(N__14460),
            .lcout(\uu2.w_data_i_0_tzZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m59_bm_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m59_bm_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m59_bm_LC_5_9_0 .LUT_INIT=16'b0000001101011111;
    LogicCell40 \Lab_UT.bcd2segment1.m59_bm_LC_5_9_0  (
            .in0(N__9612),
            .in1(N__18096),
            .in2(N__16828),
            .in3(N__16695),
            .lcout(\Lab_UT.bcd2segment1.m59_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m52_am_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m52_am_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m52_am_LC_5_9_1 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \Lab_UT.bcd2segment1.m52_am_LC_5_9_1  (
            .in0(N__16811),
            .in1(N__10446),
            .in2(N__16721),
            .in3(N__14166),
            .lcout(\Lab_UT.bcd2segment1.m52_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_0_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_0_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_0_LC_5_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.alarmchar_0_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__10584),
            .in2(_gnd_net_),
            .in3(N__10808),
            .lcout(\Lab_UT.alarmcharZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18451),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_4_LC_5_9_3 .LUT_INIT=16'b1110111110101011;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_LC_5_9_3  (
            .in0(N__10350),
            .in1(N__13329),
            .in2(N__13314),
            .in3(N__13251),
            .lcout(\Lab_UT.dictrl.state_retZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18451),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_5_9_4 .LUT_INIT=16'b1000100010001101;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_5_9_4  (
            .in0(N__9828),
            .in1(N__9873),
            .in2(N__10854),
            .in3(N__10751),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_5_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_5_9_5  (
            .in0(N__9874),
            .in1(N__9827),
            .in2(_gnd_net_),
            .in3(N__10561),
            .lcout(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ),
            .ltout(\Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_74_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_74_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_74_LC_5_9_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__G_74_LC_5_9_6  (
            .in0(N__9829),
            .in1(N__9568),
            .in2(N__9552),
            .in3(N__10349),
            .lcout(\Lab_UT.dictrl.G_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m59_am_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m59_am_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m59_am_LC_5_9_7 .LUT_INIT=16'b1011111110110000;
    LogicCell40 \Lab_UT.bcd2segment1.m59_am_LC_5_9_7  (
            .in0(N__16810),
            .in1(N__14255),
            .in2(N__16720),
            .in3(N__16311),
            .lcout(\Lab_UT.bcd2segment1.m59_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_5_10_0 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_1_LC_5_10_0  (
            .in0(N__10847),
            .in1(N__9840),
            .in2(N__9888),
            .in3(N__10752),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_5_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_0_LC_5_10_1  (
            .in0(N__9883),
            .in1(N__9838),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_5_10_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_5_10_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_LC_5_10_2  (
            .in0(N__10563),
            .in1(N__9884),
            .in2(_gnd_net_),
            .in3(N__9839),
            .lcout(\Lab_UT.dictrl.alarmstate_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.dispString.cnt_3_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_3_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_3_LC_5_10_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \Lab_UT.dispString.cnt_3_LC_5_10_3  (
            .in0(N__16816),
            .in1(N__9797),
            .in2(N__16724),
            .in3(N__10639),
            .lcout(\Lab_UT.cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.dispString.cnt_0_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_5_10_4 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_5_10_4  (
            .in0(N__9795),
            .in1(N__16711),
            .in2(N__10656),
            .in3(N__16817),
            .lcout(\Lab_UT.cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.dispString.cnt_2_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_5_10_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_5_10_5  (
            .in0(N__16710),
            .in1(N__10635),
            .in2(_gnd_net_),
            .in3(N__9796),
            .lcout(\Lab_UT.cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18444),
            .ce(),
            .sr(N__18690));
    defparam \Lab_UT.bcd2segment1.m8_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m8_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m8_LC_5_10_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m8_LC_5_10_7  (
            .in0(N__14102),
            .in1(N__14266),
            .in2(_gnd_net_),
            .in3(N__14177),
            .lcout(\Lab_UT.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_5_LC_5_11_0 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_5_11_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_5_LC_5_11_0  (
            .in0(N__9777),
            .in1(N__10721),
            .in2(_gnd_net_),
            .in3(N__10740),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu2.l_count_6_LC_5_11_1 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_5_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.l_count_6_LC_5_11_1  (
            .in0(N__10685),
            .in1(N__9753),
            .in2(_gnd_net_),
            .in3(N__9776),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \Lab_UT.dictrl.state_ret_2_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_LC_5_11_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_LC_5_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__13293),
            .in2(_gnd_net_),
            .in3(N__13272),
            .lcout(\Lab_UT.dictrl.dicRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu0.sec_clk_LC_5_11_3 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_5_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__9643),
            .in2(_gnd_net_),
            .in3(N__9726),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu2.vram_rd_clk_LC_5_11_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_5_11_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_5_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__10059),
            .in2(_gnd_net_),
            .in3(N__10039),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu2.l_count_3_LC_5_11_6 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_5_11_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu2.l_count_3_LC_5_11_6  (
            .in0(N__9968),
            .in1(N__10040),
            .in2(N__9984),
            .in3(N__10026),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu0.delay_line_1_LC_5_11_7 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_5_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10011),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18437),
            .ce(),
            .sr(N__18691));
    defparam \uu2.l_count_2_LC_5_12_1 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_5_12_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_5_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__9980),
            .in2(_gnd_net_),
            .in3(N__9967),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18432),
            .ce(),
            .sr(N__18708));
    defparam \buart.Z_rx.hh_0_LC_5_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_5_12_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9939),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18432),
            .ce(),
            .sr(N__18708));
    defparam \uu2.l_count_8_LC_5_12_7 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_5_12_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_5_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__9907),
            .in2(_gnd_net_),
            .in3(N__9924),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18432),
            .ce(),
            .sr(N__18708));
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_5_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_5_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_0_LC_5_13_0  (
            .in0(N__16606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.next_alarmstate_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18427),
            .ce(N__9852),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_5_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_14_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13358),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18425),
            .ce(),
            .sr(N__18709));
    defparam \Lab_UT.bcd2segment1.m89_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m89_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m89_LC_6_4_1 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \Lab_UT.bcd2segment1.m89_LC_6_4_1  (
            .in0(N__19072),
            .in1(N__19362),
            .in2(N__19180),
            .in3(N__19284),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_6_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_6_4_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_93_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10179),
            .in3(N__14982),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__18659));
    defparam \Lab_UT.bcd2segment1.m92_LC_6_4_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m92_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m92_LC_6_4_3 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \Lab_UT.bcd2segment1.m92_LC_6_4_3  (
            .in0(N__19073),
            .in1(N__19363),
            .in2(N__19181),
            .in3(N__19285),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_221_LC_6_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_6_4_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_221_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10176),
            .in3(N__14981),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__18659));
    defparam \uu2.mem0.ram512X8_inst_RNO_78_LC_6_4_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_78_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_78_LC_6_4_5 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_78_LC_6_4_5  (
            .in0(N__15996),
            .in1(_gnd_net_),
            .in2(N__10164),
            .in3(N__10173),
            .lcout(\uu2.mem0.N_107_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_83_LC_6_4_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_83_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_83_LC_6_4_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_83_LC_6_4_6  (
            .in0(N__10172),
            .in1(N__10160),
            .in2(_gnd_net_),
            .in3(N__15995),
            .lcout(),
            .ltout(\uu2.mem0.N_107_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_6_4_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_6_4_7 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_59_LC_6_4_7  (
            .in0(N__11952),
            .in1(N__15906),
            .in2(N__10152),
            .in3(N__10926),
            .lcout(\uu2.mem0.N_74_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_5_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_6_5_0  (
            .in0(N__14388),
            .in1(N__10148),
            .in2(N__14532),
            .in3(N__12759),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_6_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_6_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_23_LC_6_5_2  (
            .in0(N__12074),
            .in1(N__15192),
            .in2(N__14670),
            .in3(N__15713),
            .lcout(),
            .ltout(\uu2.mem0.N_130_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_3  (
            .in0(N__14526),
            .in1(N__10113),
            .in2(N__10089),
            .in3(N__14389),
            .lcout(\uu2.mem0.N_54_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_6_5_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_6_5_4 .LUT_INIT=16'b1010000000001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_33_LC_6_5_4  (
            .in0(N__11138),
            .in1(N__12475),
            .in2(N__12770),
            .in3(N__12360),
            .lcout(),
            .ltout(\uu2.mem0.N_17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_6_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_6_5_5 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_19_LC_6_5_5  (
            .in0(N__11055),
            .in1(N__14521),
            .in2(N__10263),
            .in3(N__14387),
            .lcout(\uu2.mem0.G_13_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_5_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_6_5_7  (
            .in0(N__14525),
            .in1(N__15329),
            .in2(N__10251),
            .in3(N__14390),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_6_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_6_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_50_LC_6_6_0  (
            .in0(N__12609),
            .in1(N__16104),
            .in2(N__13919),
            .in3(N__11936),
            .lcout(\uu2.mem0.G_13_0_a3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_6_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_6_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_55_LC_6_6_1  (
            .in0(N__10437),
            .in1(N__11939),
            .in2(N__10890),
            .in3(N__10200),
            .lcout(\uu2.mem0.N_74_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_6_6_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_6_6_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_66_LC_6_6_2  (
            .in0(N__11938),
            .in1(N__13811),
            .in2(N__12477),
            .in3(N__16103),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_87_LC_6_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_87_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_87_LC_6_6_3 .LUT_INIT=16'b0001001001001001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_87_LC_6_6_3  (
            .in0(N__13810),
            .in1(N__12608),
            .in2(N__16117),
            .in3(N__12840),
            .lcout(),
            .ltout(\uu2.mem0.g0_7_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_6_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_6_6_4 .LUT_INIT=16'b0000001000001111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_62_LC_6_6_4  (
            .in0(N__14732),
            .in1(N__14277),
            .in2(N__10182),
            .in3(N__10413),
            .lcout(\uu2.mem0.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_91_LC_6_6_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_91_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_91_LC_6_6_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_91_LC_6_6_5  (
            .in0(N__13989),
            .in1(N__10430),
            .in2(N__11208),
            .in3(N__12492),
            .lcout(),
            .ltout(\uu2.mem0.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_85_LC_6_6_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_85_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_85_LC_6_6_6 .LUT_INIT=16'b1000111100000111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_85_LC_6_6_6  (
            .in0(N__15330),
            .in1(N__15573),
            .in2(N__10440),
            .in3(N__10412),
            .lcout(\uu2.mem0.N_57_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_6_6_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_6_6_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_64_LC_6_6_7  (
            .in0(N__11937),
            .in1(N__12471),
            .in2(N__13827),
            .in3(N__12341),
            .lcout(\uu2.mem0.g0_i_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_77_LC_6_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_77_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_77_LC_6_7_0 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_77_LC_6_7_0  (
            .in0(N__16014),
            .in1(N__15994),
            .in2(_gnd_net_),
            .in3(N__15924),
            .lcout(\uu2.mem0.N_98_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI64LA_1_LC_6_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI64LA_1_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI64LA_1_LC_6_7_2 .LUT_INIT=16'b1000000110000001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI64LA_1_LC_6_7_2  (
            .in0(N__10429),
            .in1(N__12839),
            .in2(N__11204),
            .in3(_gnd_net_),
            .lcout(\uu2.N_1585_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m62_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m62_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m62_LC_6_7_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.bcd2segment1.m62_LC_6_7_3  (
            .in0(N__16823),
            .in1(N__19368),
            .in2(_gnd_net_),
            .in3(N__12923),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.i6_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m68_am_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m68_am_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m68_am_LC_6_7_4 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \Lab_UT.bcd2segment1.m68_am_LC_6_7_4  (
            .in0(N__16252),
            .in1(N__16694),
            .in2(N__10404),
            .in3(N__16824),
            .lcout(\Lab_UT.bcd2segment1.m68_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIV7KP6_8_LC_6_7_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIV7KP6_8_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIV7KP6_8_LC_6_7_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIV7KP6_8_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__10339),
            .in2(_gnd_net_),
            .in3(N__15428),
            .lcout(\uu2.un21_w_addr_displaying_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_39_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__15335),
            .in2(_gnd_net_),
            .in3(N__15581),
            .lcout(\uu2.mem0.N_126_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_6_7_7 .C_ON=1'b0;
    defparam \resetGen.rst_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_6_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10395),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18455),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_6_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_6_8_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_6_8_0  (
            .in0(N__14352),
            .in1(N__10310),
            .in2(N__11180),
            .in3(N__14487),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_6_8_1 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_6_8_1 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_6_8_1  (
            .in0(N__10532),
            .in1(N__14486),
            .in2(_gnd_net_),
            .in3(N__14351),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_6_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_6_8_3 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_36_LC_6_8_3  (
            .in0(N__15187),
            .in1(N__15332),
            .in2(N__14683),
            .in3(N__15582),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_8_4 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_20_LC_6_8_4  (
            .in0(N__10467),
            .in1(N__10473),
            .in2(N__10488),
            .in3(N__14736),
            .lcout(\uu2.mem0.g1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_8_5 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_35_LC_6_8_5  (
            .in0(N__12736),
            .in1(N__11168),
            .in2(_gnd_net_),
            .in3(N__12325),
            .lcout(\uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_6_8_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_6_8_6 .LUT_INIT=16'b0001001001001001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_37_LC_6_8_6  (
            .in0(N__12326),
            .in1(N__12737),
            .in2(N__11179),
            .in3(N__12476),
            .lcout(\uu2.mem0.g0_7_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_8_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_6_8_7  (
            .in0(N__15678),
            .in1(N__11172),
            .in2(N__12755),
            .in3(N__12327),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__14578),
            .sr(N__18650));
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__10583),
            .in2(_gnd_net_),
            .in3(N__10807),
            .lcout(),
            .ltout(\Lab_UT.alarmchar9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_2_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_2_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_2_LC_6_9_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.alarmchar_2_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10461),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmcharZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18441),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m47_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m47_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m47_LC_6_9_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \Lab_UT.bcd2segment1.m47_LC_6_9_2  (
            .in0(N__19173),
            .in1(N__16790),
            .in2(_gnd_net_),
            .in3(N__13049),
            .lcout(\Lab_UT.bcd2segment1.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m36_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m36_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m36_LC_6_9_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.bcd2segment1.m36_LC_6_9_4  (
            .in0(N__16812),
            .in1(N__19287),
            .in2(_gnd_net_),
            .in3(N__12985),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.i5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m42_am_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m42_am_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m42_am_LC_6_9_5 .LUT_INIT=16'b0100011100000011;
    LogicCell40 \Lab_UT.bcd2segment1.m42_am_LC_6_9_5  (
            .in0(N__16794),
            .in1(N__16719),
            .in2(N__10665),
            .in3(N__14103),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.m42_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_6_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_6_9_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__10634),
            .in2(N__10599),
            .in3(N__16626),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18441),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m52_bm_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m52_bm_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m52_bm_LC_6_9_7 .LUT_INIT=16'b0001000000011100;
    LogicCell40 \Lab_UT.bcd2segment1.m52_bm_LC_6_9_7  (
            .in0(N__16844),
            .in1(N__16718),
            .in2(N__16822),
            .in3(N__18026),
            .lcout(\Lab_UT.bcd2segment1.m52_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m47_0_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m47_0_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m47_0_LC_6_10_0 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \Lab_UT.bcd2segment1.m47_0_LC_6_10_0  (
            .in0(N__10590),
            .in1(N__13050),
            .in2(N__17760),
            .in3(N__13628),
            .lcout(\Lab_UT.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m41_0_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m41_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m41_0_LC_6_10_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m41_0_LC_6_10_1  (
            .in0(N__12913),
            .in1(N__12967),
            .in2(_gnd_net_),
            .in3(N__16373),
            .lcout(\Lab_UT.bcd2segment1.N_42_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_10_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__10770),
            .in2(_gnd_net_),
            .in3(N__10801),
            .lcout(),
            .ltout(\Lab_UT.dictrl.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_10_3 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_10_3  (
            .in0(N__10582),
            .in1(N__10846),
            .in2(N__10566),
            .in3(N__11330),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_1_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_1_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_1_LC_6_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.alarmchar_1_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__10771),
            .in2(_gnd_net_),
            .in3(N__10803),
            .lcout(\Lab_UT.alarmcharZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18435),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m49_0_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m49_0_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m49_0_LC_6_10_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \Lab_UT.bcd2segment1.m49_0_LC_6_10_5  (
            .in0(N__12912),
            .in1(N__12966),
            .in2(_gnd_net_),
            .in3(N__16374),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m54_0_LC_6_10_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m54_0_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m54_0_LC_6_10_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.bcd2segment1.m54_0_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__13627),
            .in2(N__10812),
            .in3(N__17709),
            .lcout(\Lab_UT.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_6_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_6_10_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_6_10_7  (
            .in0(N__10802),
            .in1(N__10772),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_11_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_6_11_0  (
            .in0(N__11390),
            .in1(N__11409),
            .in2(_gnd_net_),
            .in3(N__16514),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18430),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_6_11_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_6_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__10739),
            .in2(_gnd_net_),
            .in3(N__10722),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m60_0_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m60_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m60_0_LC_6_11_2 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \Lab_UT.bcd2segment1.m60_0_LC_6_11_2  (
            .in0(N__12971),
            .in1(N__16378),
            .in2(N__11574),
            .in3(N__13626),
            .lcout(),
            .ltout(\Lab_UT.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_11_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_6_11_3  (
            .in0(N__13194),
            .in1(N__13163),
            .in2(N__10668),
            .in3(N__12972),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18430),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__11389),
            .in2(_gnd_net_),
            .in3(N__16513),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18430),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_4_LC_6_12_0 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_6_12_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \resetGen.escKey_4_LC_6_12_0  (
            .in0(N__11667),
            .in1(N__11570),
            .in2(N__11742),
            .in3(N__17752),
            .lcout(\resetGen.escKeyZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI18N1_5_LC_6_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI18N1_5_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI18N1_5_LC_6_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI18N1_5_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__11495),
            .in2(_gnd_net_),
            .in3(N__11388),
            .lcout(\buart.Z_rx.ser_clk_2 ),
            .ltout(\buart.Z_rx.ser_clk_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_12_5 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_6_12_5  (
            .in0(N__11481),
            .in1(N__17094),
            .in2(N__10860),
            .in3(N__16515),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18426),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_12_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_12_7  (
            .in0(N__11361),
            .in1(N__11408),
            .in2(N__11448),
            .in3(N__11466),
            .lcout(\buart.Z_rx.ser_clk_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state16_5_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state16_5_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state16_5_LC_6_13_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.next_state16_5_LC_6_13_0  (
            .in0(N__11731),
            .in1(N__11656),
            .in2(N__11703),
            .in3(N__11528),
            .lcout(\Lab_UT.dictrl.next_state16Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_2_0_LC_6_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_2_0_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_2_0_LC_6_13_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_2_0_LC_6_13_1  (
            .in0(N__11529),
            .in1(N__11733),
            .in2(N__11666),
            .in3(N__17741),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_6_13_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_LC_6_13_2  (
            .in0(N__17703),
            .in1(N__10824),
            .in2(N__10857),
            .in3(N__11561),
            .lcout(\Lab_UT.dictrl.next_alarmstateZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_6_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_0_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__11692),
            .in2(_gnd_net_),
            .in3(N__11599),
            .lcout(\Lab_UT.dictrl.next_alarmstate4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_3_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_3_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_3_LC_6_13_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.next_state_0_sqmuxa_3_LC_6_13_4  (
            .in0(N__17702),
            .in1(N__11530),
            .in2(N__11704),
            .in3(N__11562),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_6_13_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_6_13_5  (
            .in0(N__11660),
            .in1(N__10872),
            .in2(N__10818),
            .in3(N__17742),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIHE146_2_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIHE146_2_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIHE146_2_LC_6_13_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIHE146_2_LC_6_13_6  (
            .in0(N__14947),
            .in1(N__13427),
            .in2(N__10815),
            .in3(N__11433),
            .lcout(\Lab_UT.dictrl.next_state_set ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_0_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_0_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_0_LC_6_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_sqmuxa_0_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__11732),
            .in2(_gnd_net_),
            .in3(N__11600),
            .lcout(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_0_LC_6_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_0_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_0_LC_6_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_sqmuxa_0_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__11602),
            .in2(_gnd_net_),
            .in3(N__17739),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_LC_6_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_6_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11665),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18423),
            .ce(N__17660),
            .sr(N__18710));
    defparam \buart.Z_rx.shifter_1_LC_6_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_6_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18423),
            .ce(N__17660),
            .sr(N__18710));
    defparam \buart.Z_rx.shifter_4_LC_6_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_6_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_4_LC_6_14_6  (
            .in0(N__11603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18423),
            .ce(N__17660),
            .sr(N__18710));
    defparam \buart.Z_rx.shifter_5_LC_6_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_6_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_6_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11740),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18423),
            .ce(N__17660),
            .sr(N__18710));
    defparam \Lab_UT.bcd2segment1.m99_LC_7_3_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m99_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m99_LC_7_3_0 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \Lab_UT.bcd2segment1.m99_LC_7_3_0  (
            .in0(N__19349),
            .in1(N__19283),
            .in2(N__19179),
            .in3(N__19071),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_90_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_7_3_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_90_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10863),
            .in3(N__14980),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__18663));
    defparam \Lab_UT.bcd2segment1.segmentUQ_1_4_LC_7_3_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_1_4_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_1_4_LC_7_3_2 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_1_4_LC_7_3_2  (
            .in0(N__19348),
            .in1(N__19282),
            .in2(N__19178),
            .in3(N__19070),
            .lcout(\Lab_UT.bcd2segment1.segmentUQ_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_90_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_90_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_90_LC_7_3_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_90_LC_7_3_3  (
            .in0(N__10901),
            .in1(N__15053),
            .in2(_gnd_net_),
            .in3(N__10910),
            .lcout(),
            .ltout(\uu2.mem0.N_92_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_84_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_84_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_84_LC_7_3_4 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_84_LC_7_3_4  (
            .in0(N__11954),
            .in1(N__12220),
            .in2(N__10929),
            .in3(N__11768),
            .lcout(\uu2.mem0.m73_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_218_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_7_3_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_218_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(N__10920),
            .in2(_gnd_net_),
            .in3(N__14979),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__18663));
    defparam \uu2.mem0.ram512X8_inst_RNO_88_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_88_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_88_LC_7_3_6 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_88_LC_7_3_6  (
            .in0(N__15054),
            .in1(_gnd_net_),
            .in2(N__10914),
            .in3(N__10902),
            .lcout(),
            .ltout(\uu2.mem0.N_92_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_79_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_79_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_79_LC_7_3_7 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_79_LC_7_3_7  (
            .in0(N__11769),
            .in1(N__12222),
            .in2(N__10893),
            .in3(N__11955),
            .lcout(\uu2.mem0.m73_ns_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m26_0_LC_7_4_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m26_0_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m26_0_LC_7_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m26_0_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(N__14057),
            .in2(_gnd_net_),
            .in3(N__14243),
            .lcout(\Lab_UT.N_27_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_7_4_3 .LUT_INIT=16'b1111011010010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_40_LC_7_4_3  (
            .in0(N__15677),
            .in1(N__11163),
            .in2(N__11972),
            .in3(N__10878),
            .lcout(\uu2.mem0.i14_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_4_6 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_7_4_6  (
            .in0(N__16302),
            .in1(N__14058),
            .in2(N__13113),
            .in3(N__14244),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18491),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m106_LC_7_4_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m106_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m106_LC_7_4_7 .LUT_INIT=16'b1110110011000011;
    LogicCell40 \Lab_UT.bcd2segment1.m106_LC_7_4_7  (
            .in0(N__14242),
            .in1(N__14154),
            .in2(N__14083),
            .in3(N__16241),
            .lcout(\Lab_UT.bcd2segment1.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_7_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_7_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_34_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__15328),
            .in2(_gnd_net_),
            .in3(N__15580),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_7_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_7_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_7_5_1  (
            .in0(N__14386),
            .in1(N__14520),
            .in2(_gnd_net_),
            .in3(N__11049),
            .lcout(\uu2.mem0.N_93_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_5_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_60_LC_7_5_3  (
            .in0(N__12433),
            .in1(N__12359),
            .in2(N__13920),
            .in3(N__13826),
            .lcout(\uu2.mem0.N_67_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_7_5_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_61_LC_7_5_4  (
            .in0(N__14519),
            .in1(N__14385),
            .in2(_gnd_net_),
            .in3(N__11019),
            .lcout(),
            .ltout(\uu2.mem0.g0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_7_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_7_5_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_41_LC_7_5_5  (
            .in0(N__13932),
            .in1(N__11013),
            .in2(N__11007),
            .in3(N__11004),
            .lcout(),
            .ltout(\uu2.mem0.g0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_7_5_6 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_21_LC_7_5_6  (
            .in0(N__10998),
            .in1(N__10992),
            .in2(N__10980),
            .in3(N__12000),
            .lcout(),
            .ltout(\uu2.mem0.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_7_5_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_7_5_7  (
            .in0(N__10977),
            .in1(N__12021),
            .in2(N__10971),
            .in3(N__14289),
            .lcout(\uu2.mem0.N_66_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_7_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_7_6_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_42_LC_7_6_0  (
            .in0(N__10956),
            .in1(N__15331),
            .in2(N__10938),
            .in3(N__15577),
            .lcout(\uu2.mem0.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_7_6_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_7_6_1 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_65_LC_7_6_1  (
            .in0(N__12331),
            .in1(N__13904),
            .in2(_gnd_net_),
            .in3(N__13816),
            .lcout(\uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_RNINBDH1_LC_7_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNINBDH1_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNINBDH1_LC_7_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNINBDH1_LC_7_6_2  (
            .in0(N__11130),
            .in1(N__12426),
            .in2(N__13917),
            .in3(N__12330),
            .lcout(\uu2.N_67_1_0 ),
            .ltout(\uu2.N_67_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_7_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_7_6_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_25_LC_7_6_3  (
            .in0(N__15651),
            .in1(_gnd_net_),
            .in2(N__11076),
            .in3(N__11064),
            .lcout(\uu2.mem0.N_55_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_7_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_7_6_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_48_LC_7_6_4  (
            .in0(N__13900),
            .in1(N__12425),
            .in2(_gnd_net_),
            .in3(N__12329),
            .lcout(\uu2.mem0.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_LC_7_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_7_6_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_displaying_1_LC_7_6_5  (
            .in0(N__15652),
            .in1(N__11131),
            .in2(_gnd_net_),
            .in3(N__15451),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__18657));
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_6_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_LC_7_6_6  (
            .in0(N__15452),
            .in1(_gnd_net_),
            .in2(N__13828),
            .in3(N__15653),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__18657));
    defparam \uu2.w_addr_displaying_1_rep1_RNIKGI51_LC_7_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIKGI51_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIKGI51_LC_7_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIKGI51_LC_7_6_7  (
            .in0(N__12424),
            .in1(N__16102),
            .in2(N__13918),
            .in3(N__13815),
            .lcout(\uu2.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m118_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m118_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m118_LC_7_7_0 .LUT_INIT=16'b1110110111001010;
    LogicCell40 \Lab_UT.bcd2segment1.m118_LC_7_7_0  (
            .in0(N__14245),
            .in1(N__14161),
            .in2(N__14098),
            .in3(N__16242),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_250_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_7_7_1 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_7_7_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_296_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11058),
            .in3(N__14935),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__18656));
    defparam \Lab_UT.bcd2segment1.m97_0_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m97_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m97_0_LC_7_7_2 .LUT_INIT=16'b0000100110000010;
    LogicCell40 \Lab_UT.bcd2segment1.m97_0_LC_7_7_2  (
            .in0(N__14246),
            .in1(N__14162),
            .in2(N__14099),
            .in3(N__16243),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_7_7_3 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_7_7_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_40_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11244),
            .in3(N__14936),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__18656));
    defparam \uu2.mem0.ram512X8_inst_RNO_74_LC_7_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_74_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_74_LC_7_7_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_74_LC_7_7_4  (
            .in0(N__11237),
            .in1(_gnd_net_),
            .in2(N__11226),
            .in3(N__14784),
            .lcout(\uu2.mem0.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIJVK41_40_LC_7_7_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJVK41_40_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJVK41_40_LC_7_7_5 .LUT_INIT=16'b0001001111010011;
    LogicCell40 \uu2.bitmap_RNIJVK41_40_LC_7_7_5  (
            .in0(N__11241),
            .in1(N__13217),
            .in2(N__12221),
            .in3(N__11222),
            .lcout(),
            .ltout(\uu2.m95_i_m2_i_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI19S42_34_LC_7_7_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI19S42_34_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI19S42_34_LC_7_7_6 .LUT_INIT=16'b1111000000110101;
    LogicCell40 \uu2.bitmap_RNI19S42_34_LC_7_7_6  (
            .in0(N__12525),
            .in1(N__12549),
            .in2(N__11214),
            .in3(N__12213),
            .lcout(\uu2.N_16 ),
            .ltout(\uu2.N_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_7_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_7_7_7 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_57_LC_7_7_7  (
            .in0(N__15183),
            .in1(N__12432),
            .in2(N__11211),
            .in3(N__11993),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_7_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_7_8_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_LC_7_8_0  (
            .in0(N__15679),
            .in1(N__12731),
            .in2(N__11181),
            .in3(N__12214),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .ce(N__14579),
            .sr(N__18651));
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_7_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_7_8_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_3_LC_7_8_1  (
            .in0(N__11151),
            .in1(N__15681),
            .in2(N__12753),
            .in3(N__11203),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .ce(N__14579),
            .sr(N__18651));
    defparam \uu2.w_addr_displaying_3_rep2_nesr_LC_7_8_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep2_nesr_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep2_nesr_LC_7_8_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_3_rep2_nesr_LC_7_8_2  (
            .in0(N__15680),
            .in1(N__11152),
            .in2(N__16116),
            .in3(N__12732),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .ce(N__14579),
            .sr(N__18651));
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_7_8_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_7_8_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_nesr_LC_7_8_3  (
            .in0(N__15333),
            .in1(N__15189),
            .in2(N__15399),
            .in3(N__14786),
            .lcout(\uu2.w_addr_displaying_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .ce(N__14579),
            .sr(N__18651));
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_7_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_7_8_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_8_LC_7_8_4  (
            .in0(N__15188),
            .in1(N__15334),
            .in2(N__13221),
            .in3(N__15396),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1_nesrC_net ),
            .ce(N__14579),
            .sr(N__18651));
    defparam CONSTANT_ONE_LUT4_LC_7_8_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_8_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_7_9_0 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_0_LC_7_9_0  (
            .in0(N__18091),
            .in1(N__18025),
            .in2(N__18178),
            .in3(N__19436),
            .lcout(\Lab_UT.bcd2segment2.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_7_9_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_7_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_70_LC_7_9_1  (
            .in0(N__14793),
            .in1(N__12651),
            .in2(_gnd_net_),
            .in3(N__13233),
            .lcout(\uu2.mem0.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_7_9_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_7_9_2  (
            .in0(N__13102),
            .in1(N__11297),
            .in2(N__16295),
            .in3(N__16254),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18452),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_7_9_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_7_9_3  (
            .in0(N__16167),
            .in1(N__14160),
            .in2(N__11301),
            .in3(N__13098),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18452),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_7_9_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_7_9_4  (
            .in0(N__16288),
            .in1(_gnd_net_),
            .in2(N__13106),
            .in3(N__14241),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18452),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.un1_num_1_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.un1_num_1_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.un1_num_1_LC_7_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.bcd2segment2.un1_num_1_LC_7_9_5  (
            .in0(N__19435),
            .in1(N__18090),
            .in2(N__18027),
            .in3(N__18166),
            .lcout(\Lab_UT.zero ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_71_LC_7_9_6  (
            .in0(N__14785),
            .in1(N__12524),
            .in2(_gnd_net_),
            .in3(N__12548),
            .lcout(\uu2.mem0.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_7_9_7 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_7_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.escKey_LC_7_9_7  (
            .in0(N__11757),
            .in1(N__11283),
            .in2(_gnd_net_),
            .in3(N__17058),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_7_10_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_7_10_0 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_67_LC_7_10_0  (
            .in0(N__13913),
            .in1(N__16108),
            .in2(_gnd_net_),
            .in3(N__13829),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNIASM81_2_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNIASM81_2_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNIASM81_2_LC_7_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNIASM81_2_LC_7_10_1  (
            .in0(N__12959),
            .in1(N__16360),
            .in2(N__12901),
            .in3(N__14216),
            .lcout(),
            .ltout(\Lab_UT.didp.did_alarmMatch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIUG9D3_1_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIUG9D3_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIUG9D3_1_LC_7_10_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIUG9D3_1_LC_7_10_2  (
            .in0(N__14076),
            .in1(N__11322),
            .in2(N__11340),
            .in3(N__11337),
            .lcout(\Lab_UT.alarmMatch ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNISKK51_3_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNISKK51_3_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNISKK51_3_LC_7_10_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNISKK51_3_LC_7_10_3  (
            .in0(N__13051),
            .in1(N__14136),
            .in2(_gnd_net_),
            .in3(N__16214),
            .lcout(\Lab_UT.didp.countrce3.did_alarmMatch_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_7_10_4  (
            .in0(N__11316),
            .in1(N__13162),
            .in2(N__13190),
            .in3(N__13052),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18445),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m65_0_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m65_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m65_0_LC_7_10_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.bcd2segment1.m65_0_LC_7_10_5  (
            .in0(N__13629),
            .in1(N__16361),
            .in2(_gnd_net_),
            .in3(N__11532),
            .lcout(),
            .ltout(\Lab_UT.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_10_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_7_10_6  (
            .in0(N__16362),
            .in1(N__13182),
            .in2(N__11310),
            .in3(N__13158),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18445),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_10_7 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_7_10_7  (
            .in0(N__12883),
            .in1(N__13183),
            .in2(N__13164),
            .in3(N__11307),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18445),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_7_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__17877),
            .in2(_gnd_net_),
            .in3(N__18746),
            .lcout(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI72HD1_1_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI72HD1_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI72HD1_1_LC_7_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI72HD1_1_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__11421),
            .in2(_gnd_net_),
            .in3(N__17948),
            .lcout(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_7_11_2 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_1_LC_7_11_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_7_11_2  (
            .in0(N__17949),
            .in1(N__17547),
            .in2(N__11424),
            .in3(N__17804),
            .lcout(\Lab_UT.dictrl.next_state_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18438),
            .ce(N__17494),
            .sr(N__13647));
    defparam \Lab_UT.dictrl.state_0_RNITK4F_1_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNITK4F_1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNITK4F_1_LC_7_11_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNITK4F_1_LC_7_11_3  (
            .in0(N__16907),
            .in1(N__13776),
            .in2(_gnd_net_),
            .in3(N__13507),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_RNIS90D1_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNIS90D1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNIS90D1_LC_7_11_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNIS90D1_LC_7_11_4  (
            .in0(N__18908),
            .in1(N__16908),
            .in2(N__11415),
            .in3(N__18953),
            .lcout(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1 ),
            .ltout(\Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIR0FR1_3_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIR0FR1_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIR0FR1_3_LC_7_11_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIR0FR1_3_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11412),
            .in3(N__16551),
            .lcout(\Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_7_11_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_7_11_6  (
            .in0(N__18983),
            .in1(N__18952),
            .in2(_gnd_net_),
            .in3(N__18877),
            .lcout(\Lab_UT.Run ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_7_12_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__11407),
            .in2(N__11391),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_7_12_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_7_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__11465),
            .in2(_gnd_net_),
            .in3(N__11364),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_2  (
            .in0(N__16487),
            .in1(N__11357),
            .in2(_gnd_net_),
            .in3(N__11346),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__18433),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_12_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__11447),
            .in2(_gnd_net_),
            .in3(N__11343),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__11496),
            .in2(_gnd_net_),
            .in3(N__11484),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_7_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_7_12_5 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_7_12_5  (
            .in0(N__16485),
            .in1(N__17087),
            .in2(N__11475),
            .in3(N__17121),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18433),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIPU6T9_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIPU6T9_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIPU6T9_LC_7_12_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIPU6T9_LC_7_12_6  (
            .in0(N__17945),
            .in1(N__17911),
            .in2(N__17870),
            .in3(N__17796),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_7 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_7  (
            .in0(N__16486),
            .in1(N__17122),
            .in2(N__17100),
            .in3(N__11454),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18433),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_LC_7_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_7_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_7_LC_7_13_0  (
            .in0(N__13377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18428),
            .ce(N__17653),
            .sr(N__18711));
    defparam \buart.Z_rx.shifter_6_LC_7_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_7_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_6_LC_7_13_1  (
            .in0(N__11702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18428),
            .ce(N__17653),
            .sr(N__18711));
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_7_13_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \Lab_UT.dictrl.state_0_RNILGF17_3_LC_7_13_3  (
            .in0(N__13640),
            .in1(N__11748),
            .in2(N__14934),
            .in3(N__11621),
            .lcout(\Lab_UT.dictrl.next_state_set_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_13_5 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_13_5  (
            .in0(N__13586),
            .in1(N__13770),
            .in2(_gnd_net_),
            .in3(N__13565),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxa_1 ),
            .ltout(\Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIJ9317_2_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIJ9317_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIJ9317_2_LC_7_13_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIJ9317_2_LC_7_13_6  (
            .in0(N__11622),
            .in1(N__14886),
            .in2(N__11427),
            .in3(N__17465),
            .lcout(\Lab_UT.dictrl.next_state_set_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_5_LC_7_13_7 .C_ON=1'b0;
    defparam \resetGen.escKey_5_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_5_LC_7_13_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \resetGen.escKey_5_LC_7_13_7  (
            .in0(N__17704),
            .in1(N__11531),
            .in2(N__11706),
            .in3(N__11610),
            .lcout(\resetGen.escKeyZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNICJTA2_3_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNICJTA2_3_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNICJTA2_3_LC_7_14_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_RNICJTA2_3_LC_7_14_0  (
            .in0(N__13548),
            .in1(N__13585),
            .in2(_gnd_net_),
            .in3(N__13564),
            .lcout(\Lab_UT.dictrl.next_state_set_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_4_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_4_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_4_LC_7_14_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_sqmuxa_4_LC_7_14_1  (
            .in0(N__11741),
            .in1(N__11524),
            .in2(N__11705),
            .in3(N__11560),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_5_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_5_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_5_LC_7_14_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_sqmuxa_5_LC_7_14_2  (
            .in0(N__11661),
            .in1(N__11631),
            .in2(N__11625),
            .in3(N__17686),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNI0MRT_1_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNI0MRT_1_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNI0MRT_1_LC_7_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNI0MRT_1_LC_7_14_5  (
            .in0(N__18969),
            .in1(N__16905),
            .in2(_gnd_net_),
            .in3(N__13516),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_state_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIS90D1_2_LC_7_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIS90D1_2_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIS90D1_2_LC_7_14_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIS90D1_2_LC_7_14_6  (
            .in0(N__13771),
            .in1(N__16906),
            .in2(N__11613),
            .in3(N__18904),
            .lcout(\Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state16_4_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state16_4_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state16_4_LC_7_14_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state16_4_LC_7_14_7  (
            .in0(N__11601),
            .in1(N__11559),
            .in2(N__17701),
            .in3(N__17740),
            .lcout(\Lab_UT.dictrl.next_state16Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_7_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11569),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18424),
            .ce(N__17661),
            .sr(N__18712));
    defparam \Lab_UT.bcd2segment1.m84_0_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m84_0_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m84_0_LC_8_3_0 .LUT_INIT=16'b0001010101100110;
    LogicCell40 \Lab_UT.bcd2segment1.m84_0_LC_8_3_0  (
            .in0(N__13063),
            .in1(N__12920),
            .in2(N__16408),
            .in3(N__13000),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_127_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_8_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_8_3_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_162_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11790),
            .in3(N__14989),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_162C_net ),
            .ce(),
            .sr(N__18666));
    defparam \Lab_UT.bcd2segment1.m87_0_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m87_0_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m87_0_LC_8_3_2 .LUT_INIT=16'b0000010001100111;
    LogicCell40 \Lab_UT.bcd2segment1.m87_0_LC_8_3_2  (
            .in0(N__13064),
            .in1(N__12921),
            .in2(N__16409),
            .in3(N__13001),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_66_LC_8_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_8_3_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_66_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11787),
            .in3(N__14991),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_162C_net ),
            .ce(),
            .sr(N__18666));
    defparam \Lab_UT.bcd2segment1.m90_0_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m90_0_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m90_0_LC_8_3_4 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \Lab_UT.bcd2segment1.m90_0_LC_8_3_4  (
            .in0(N__13065),
            .in1(N__12922),
            .in2(N__16410),
            .in3(N__13002),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_194_LC_8_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_8_3_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_194_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11784),
            .in3(N__14990),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_162C_net ),
            .ce(),
            .sr(N__18666));
    defparam \uu2.bitmap_RNIIGUI_66_LC_8_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIIGUI_66_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIIGUI_66_LC_8_3_6 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \uu2.bitmap_RNIIGUI_66_LC_8_3_6  (
            .in0(N__11781),
            .in1(N__15044),
            .in2(_gnd_net_),
            .in3(N__11775),
            .lcout(\uu2.N_101_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m93_0_LC_8_3_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m93_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m93_0_LC_8_3_7 .LUT_INIT=16'b0000000101101011;
    LogicCell40 \Lab_UT.bcd2segment1.m93_0_LC_8_3_7  (
            .in0(N__12999),
            .in1(N__16398),
            .in2(N__12924),
            .in3(N__13062),
            .lcout(\Lab_UT.bcd2segment1.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m101_LC_8_4_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m101_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m101_LC_8_4_0 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \Lab_UT.bcd2segment1.m101_LC_8_4_0  (
            .in0(N__14259),
            .in1(N__14180),
            .in2(N__14084),
            .in3(N__16255),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_8_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_8_4_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_75_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11760),
            .in3(N__14985),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_75C_net ),
            .ce(),
            .sr(N__18664));
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_8_4_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_8_4_2 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \Lab_UT.bcd2segment3.segment_0_2_LC_8_4_2  (
            .in0(N__14260),
            .in1(N__14181),
            .in2(N__14085),
            .in3(N__16256),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_203_LC_8_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_8_4_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_203_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11982),
            .in3(N__14983),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_75C_net ),
            .ce(),
            .sr(N__18664));
    defparam \uu2.bitmap_RNIC6T81_212_LC_8_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIC6T81_212_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIC6T81_212_LC_8_4_4 .LUT_INIT=16'b1101110100000011;
    LogicCell40 \uu2.bitmap_RNIC6T81_212_LC_8_4_4  (
            .in0(N__11874),
            .in1(N__15992),
            .in2(N__12663),
            .in3(N__13701),
            .lcout(),
            .ltout(\uu2.N_1580_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIL4F73_3_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIL4F73_3_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIL4F73_3_LC_8_4_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIL4F73_3_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__12368),
            .in2(N__11979),
            .in3(N__11880),
            .lcout(\uu2.N_77_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIPIHG1_75_LC_8_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_8_4_6 .LUT_INIT=16'b0101111100100010;
    LogicCell40 \uu2.bitmap_RNIPIHG1_75_LC_8_4_6  (
            .in0(N__11953),
            .in1(N__11895),
            .in2(N__11889),
            .in3(N__13995),
            .lcout(\uu2.N_1581_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_212_LC_8_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_8_4_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \uu2.bitmap_212_LC_8_4_7  (
            .in0(N__18195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14984),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_75C_net ),
            .ce(),
            .sr(N__18664));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_8_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_8_5_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_8_5_0  (
            .in0(N__15157),
            .in1(N__12064),
            .in2(N__14669),
            .in3(N__11796),
            .lcout(),
            .ltout(\uu2.mem0.N_134_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_8_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_8_5_1 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__11868),
            .in2(N__11847),
            .in3(N__11843),
            .lcout(\uu2.mem0.N_60_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_5_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_28_LC_8_5_2  (
            .in0(N__15675),
            .in1(N__12257),
            .in2(_gnd_net_),
            .in3(N__15711),
            .lcout(\uu2.mem0.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIF00Q_5_LC_8_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIF00Q_5_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIF00Q_5_LC_8_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIF00Q_5_LC_8_5_3  (
            .in0(N__15273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15550),
            .lcout(\uu2.N_126 ),
            .ltout(\uu2.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_5_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_5_4 .LUT_INIT=16'b0000000001110110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_46_LC_8_5_4  (
            .in0(N__15156),
            .in1(N__14652),
            .in2(N__12153),
            .in3(N__15712),
            .lcout(\uu2.mem0.bitmap_pmux_u_i_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_5_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_8_5_5  (
            .in0(N__14531),
            .in1(N__15676),
            .in2(N__14397),
            .in3(N__12150),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_8_5_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_8_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_44_LC_8_5_6  (
            .in0(N__12099),
            .in1(N__12087),
            .in2(_gnd_net_),
            .in3(N__12063),
            .lcout(),
            .ltout(\uu2.mem0.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_8_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_8_5_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_24_LC_8_5_7  (
            .in0(N__14697),
            .in1(N__12045),
            .in2(N__12030),
            .in3(N__12027),
            .lcout(\uu2.mem0.g0_7_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_8_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_8_6_0 .LUT_INIT=16'b1110101011101111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_58_LC_8_6_0  (
            .in0(N__12428),
            .in1(N__11994),
            .in2(N__15190),
            .in3(N__12015),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_8_6_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_8_6_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_38_LC_8_6_1  (
            .in0(N__16047),
            .in1(_gnd_net_),
            .in2(N__12009),
            .in3(N__12006),
            .lcout(\uu2.mem0.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI43641_162_LC_8_6_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI43641_162_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI43641_162_LC_8_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNI43641_162_LC_8_6_2  (
            .in0(N__12216),
            .in1(N__13676),
            .in2(_gnd_net_),
            .in3(N__12245),
            .lcout(\uu2.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_73_LC_8_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_73_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_73_LC_8_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_73_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__12594),
            .in2(_gnd_net_),
            .in3(N__12215),
            .lcout(\uu2.mem0.m317_0_a6_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_LC_8_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_rep1_LC_8_6_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_LC_8_6_4  (
            .in0(N__12595),
            .in1(N__12772),
            .in2(N__12367),
            .in3(N__12512),
            .lcout(\uu2.w_addr_displaying_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__18660));
    defparam \uu2.w_addr_displaying_4_LC_8_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_8_6_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_4_LC_8_6_5  (
            .in0(N__12447),
            .in1(N__12354),
            .in2(N__12777),
            .in3(N__12511),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__18660));
    defparam \uu2.w_addr_displaying_fast_4_LC_8_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_4_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_4_LC_8_6_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_4_LC_8_6_6  (
            .in0(N__12358),
            .in1(N__12776),
            .in2(N__12513),
            .in3(N__12491),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__18660));
    defparam \uu2.w_addr_displaying_2_rep1_RNI01H61_LC_8_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNI01H61_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNI01H61_LC_8_6_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNI01H61_LC_8_6_7  (
            .in0(N__13912),
            .in1(N__12427),
            .in2(_gnd_net_),
            .in3(N__12353),
            .lcout(\uu2.N_9_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_75_LC_8_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_75_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_75_LC_8_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_75_LC_8_7_0  (
            .in0(N__12208),
            .in1(N__13677),
            .in2(_gnd_net_),
            .in3(N__12246),
            .lcout(),
            .ltout(\uu2.mem0.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_8_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_8_7_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_54_LC_8_7_1  (
            .in0(N__15124),
            .in1(N__12228),
            .in2(N__12231),
            .in3(N__12601),
            .lcout(\uu2.mem0.m317_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_76_LC_8_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_76_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_76_LC_8_7_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_76_LC_8_7_2  (
            .in0(N__12207),
            .in1(N__15973),
            .in2(N__12607),
            .in3(N__16041),
            .lcout(\uu2.mem0.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_72_LC_8_7_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_72_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_72_LC_8_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_72_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__15966),
            .in2(_gnd_net_),
            .in3(N__12209),
            .lcout(),
            .ltout(\uu2.mem0.m317_0_a6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_7_4 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_51_LC_8_7_4  (
            .in0(N__12599),
            .in1(N__12162),
            .in2(N__12639),
            .in3(N__12636),
            .lcout(),
            .ltout(\uu2.mem0.N_11_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_29_LC_8_7_5  (
            .in0(N__12627),
            .in1(N__15003),
            .in2(N__12621),
            .in3(N__12564),
            .lcout(\uu2.mem0.N_6_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_7_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_53_LC_8_7_6  (
            .in0(N__12600),
            .in1(N__16115),
            .in2(N__15158),
            .in3(N__12570),
            .lcout(\uu2.mem0.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_31_LC_8_7_7  (
            .in0(N__15313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15560),
            .lcout(\uu2.mem0.g1_2_2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_34_LC_8_8_0 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_8_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_34_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__13083),
            .in2(_gnd_net_),
            .in3(N__14951),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.bitmap_69_LC_8_8_1 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_8_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_69_LC_8_8_1  (
            .in0(N__14952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13074),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.bitmap_197_LC_8_8_2 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_8_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_197_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__12849),
            .in2(_gnd_net_),
            .in3(N__14948),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.bitmap_290_LC_8_8_3 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_8_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_290_LC_8_8_3  (
            .in0(N__14949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12537),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.bitmap_308_LC_8_8_4 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_8_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_308_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__17574),
            .in2(_gnd_net_),
            .in3(N__14950),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.w_addr_displaying_2_rep1_LC_8_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_rep1_LC_8_8_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_LC_8_8_5  (
            .in0(N__12808),
            .in1(N__13887),
            .in2(_gnd_net_),
            .in3(N__15472),
            .lcout(\uu2.w_addr_displaying_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.w_addr_displaying_fast_2_LC_8_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_8_8_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_8_8_6  (
            .in0(N__15473),
            .in1(N__12809),
            .in2(_gnd_net_),
            .in3(N__12832),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \uu2.w_addr_displaying_2_LC_8_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_8_8_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_displaying_2_LC_8_8_7  (
            .in0(N__12807),
            .in1(N__12727),
            .in2(_gnd_net_),
            .in3(N__15471),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__18654));
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_8_9_0 .LUT_INIT=16'b1110100111100001;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_6_LC_8_9_0  (
            .in0(N__19432),
            .in1(N__18171),
            .in2(N__18021),
            .in3(N__18089),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_180_LC_8_9_1 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_8_9_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_180_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12675),
            .in3(N__14900),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_180C_net ),
            .ce(),
            .sr(N__18658));
    defparam \uu2.bitmap_52_LC_8_9_3 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_8_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_52_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__12672),
            .in2(_gnd_net_),
            .in3(N__14902),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_180C_net ),
            .ce(),
            .sr(N__18658));
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_8_9_4 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_1_LC_8_9_4  (
            .in0(N__19431),
            .in1(N__18170),
            .in2(N__18020),
            .in3(N__18087),
            .lcout(\Lab_UT.bcd2segment2.segment_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_8_9_5 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_2_LC_8_9_5  (
            .in0(N__18088),
            .in1(N__18003),
            .in2(N__18179),
            .in3(N__19433),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_8_9_6 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_8_9_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.bitmap_215_LC_8_9_6  (
            .in0(N__14901),
            .in1(_gnd_net_),
            .in2(N__12666),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_180C_net ),
            .ce(),
            .sr(N__18658));
    defparam \uu2.mem0.ram512X8_inst_RNO_89_LC_8_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_89_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_89_LC_8_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_89_LC_8_9_7  (
            .in0(N__12650),
            .in1(N__13232),
            .in2(_gnd_net_),
            .in3(N__13216),
            .lcout(\uu2.mem0.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m39_e_2_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m39_e_2_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m39_e_2_LC_8_10_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.bcd2segment1.m39_e_2_LC_8_10_0  (
            .in0(N__13048),
            .in1(N__16229),
            .in2(N__16387),
            .in3(N__18743),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m39_e_3_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m39_e_3_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m39_e_3_LC_8_10_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \Lab_UT.bcd2segment1.m39_e_3_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__12889),
            .in2(N__13200),
            .in3(N__12989),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_3_LC_8_10_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_8_10_2  (
            .in0(N__13130),
            .in1(N__18777),
            .in2(N__13197),
            .in3(N__18745),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18453),
            .ce(),
            .sr(N__18223));
    defparam \Lab_UT.didp.ce_3_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_8_10_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_8_10_3  (
            .in0(N__16230),
            .in1(N__13126),
            .in2(_gnd_net_),
            .in3(N__18776),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18453),
            .ce(),
            .sr(N__18223));
    defparam \Lab_UT.didp.reset_2_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_2_LC_8_10_4 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_8_10_4  (
            .in0(N__18775),
            .in1(N__16231),
            .in2(N__13131),
            .in3(N__18744),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18453),
            .ce(),
            .sr(N__18223));
    defparam \Lab_UT.bcd2segment1.m76_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m76_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m76_LC_8_10_5 .LUT_INIT=16'b0010000110010000;
    LogicCell40 \Lab_UT.bcd2segment1.m76_LC_8_10_5  (
            .in0(N__13043),
            .in1(N__12987),
            .in2(N__16382),
            .in3(N__12887),
            .lcout(\Lab_UT.bcd2segment1.N_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m76_0_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m76_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m76_0_LC_8_10_6 .LUT_INIT=16'b0100011110011111;
    LogicCell40 \Lab_UT.bcd2segment1.m76_0_LC_8_10_6  (
            .in0(N__12986),
            .in1(N__16363),
            .in2(N__12902),
            .in3(N__13042),
            .lcout(\Lab_UT.bcd2segment1.N_229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m81_0_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m81_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m81_0_LC_8_10_7 .LUT_INIT=16'b0111010111111011;
    LogicCell40 \Lab_UT.bcd2segment1.m81_0_LC_8_10_7  (
            .in0(N__13044),
            .in1(N__12988),
            .in2(N__16383),
            .in3(N__12888),
            .lcout(\Lab_UT.bcd2segment1.N_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_8_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__13239),
            .in2(_gnd_net_),
            .in3(N__13408),
            .lcout(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ),
            .ltout(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIQ35U8_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIQ35U8_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIQ35U8_LC_8_11_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIQ35U8_LC_8_11_2  (
            .in0(N__13409),
            .in1(N__17874),
            .in2(N__13332),
            .in3(N__13456),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_0 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIFPRO41_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIFPRO41_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIFPRO41_LC_8_11_3 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIFPRO41_LC_8_11_3  (
            .in0(N__13265),
            .in1(N__13292),
            .in2(N__13317),
            .in3(N__13304),
            .lcout(\Lab_UT.dictrl.un1_state_21_reti_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIQCSRA_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIQCSRA_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIQCSRA_LC_8_11_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIQCSRA_LC_8_11_4  (
            .in0(N__17340),
            .in1(N__17875),
            .in2(N__17305),
            .in3(N__17525),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNI2AJ17_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNI2AJ17_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNI2AJ17_LC_8_11_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNI2AJ17_LC_8_11_5  (
            .in0(N__16998),
            .in1(N__16959),
            .in2(N__17886),
            .in3(N__16936),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_3 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIR8QUG_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIR8QUG_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIR8QUG_LC_8_11_6 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIR8QUG_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13275),
            .in3(N__13264),
            .lcout(\Lab_UT.dictrl.dicRun_2_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_8_11_7 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_0_LC_8_11_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_8_11_7  (
            .in0(N__13457),
            .in1(N__17548),
            .in2(N__13475),
            .in3(N__13410),
            .lcout(\Lab_UT.dictrl.next_state_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18446),
            .ce(N__17493),
            .sr(N__13428));
    defparam \Lab_UT.dictrl.state_0_1_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_LC_8_12_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_LC_8_12_1  (
            .in0(N__17946),
            .in1(N__17912),
            .in2(N__17876),
            .in3(N__17803),
            .lcout(\Lab_UT.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18439),
            .ce(),
            .sr(N__18694));
    defparam \Lab_UT.dictrl.state_0_3_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_LC_8_12_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_LC_8_12_2  (
            .in0(N__17002),
            .in1(N__16937),
            .in2(N__16977),
            .in3(N__17861),
            .lcout(\Lab_UT.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18439),
            .ce(),
            .sr(N__18694));
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_12_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_12_4 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_8_12_4  (
            .in0(N__17521),
            .in1(N__17859),
            .in2(N__17306),
            .in3(N__17339),
            .lcout(\Lab_UT.state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18439),
            .ce(),
            .sr(N__18694));
    defparam \Lab_UT.dictrl.state_0_0_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_LC_8_12_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_LC_8_12_5  (
            .in0(N__17860),
            .in1(N__13407),
            .in2(N__13476),
            .in3(N__13458),
            .lcout(\Lab_UT.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18439),
            .ce(),
            .sr(N__18694));
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_8_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_8_12_6 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_3_LC_8_12_6  (
            .in0(N__17410),
            .in1(N__17368),
            .in2(N__16149),
            .in3(N__16483),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_3_LC_8_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_3_LC_8_12_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_3_LC_8_12_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \buart.Z_rx.bitcount_3_LC_8_12_7  (
            .in0(N__16484),
            .in1(N__17021),
            .in2(N__13431),
            .in3(N__17411),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18439),
            .ce(),
            .sr(N__18694));
    defparam \Lab_UT.bcd2segment1.m72_0_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m72_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m72_0_LC_8_13_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.bcd2segment1.m72_0_LC_8_13_0  (
            .in0(N__18894),
            .in1(N__13505),
            .in2(N__13389),
            .in3(N__16878),
            .lcout(\Lab_UT.m72_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIDH8U_1_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIDH8U_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIDH8U_1_LC_8_13_1 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIDH8U_1_LC_8_13_1  (
            .in0(N__13506),
            .in1(N__18955),
            .in2(N__16893),
            .in3(N__18896),
            .lcout(\Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m29_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m29_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m29_LC_8_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.bcd2segment1.m29_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__13531),
            .in2(_gnd_net_),
            .in3(N__13766),
            .lcout(\Lab_UT.un1_state_13 ),
            .ltout(\Lab_UT.un1_state_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_RNIAD2V_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_RNIAD2V_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_RNIAD2V_LC_8_13_3 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_RNIAD2V_LC_8_13_3  (
            .in0(N__17773),
            .in1(N__18893),
            .in2(N__13380),
            .in3(N__13338),
            .lcout(\Lab_UT.dictrl.state_ret_1_RNIAD2VZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_8_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_8_13_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.hh_RNI065O1_0_LC_8_13_5  (
            .in0(N__13376),
            .in1(N__13359),
            .in2(_gnd_net_),
            .in3(N__17139),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIENNE_1_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIENNE_1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIENNE_1_LC_8_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIENNE_1_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__13504),
            .in2(_gnd_net_),
            .in3(N__16877),
            .lcout(\Lab_UT.dictrl.un1_state_11 ),
            .ltout(\Lab_UT.dictrl.un1_state_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_RNITFCD1_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_RNITFCD1_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_RNITFCD1_LC_8_13_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_RNITFCD1_LC_8_13_7  (
            .in0(N__17774),
            .in1(N__18954),
            .in2(N__13650),
            .in3(N__18895),
            .lcout(\Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m47_e_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m47_e_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m47_e_LC_8_14_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m47_e_LC_8_14_0  (
            .in0(N__18903),
            .in1(N__17775),
            .in2(N__13772),
            .in3(N__16884),
            .lcout(\Lab_UT.bcd2segment1.N_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m68_0_ns_1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m68_0_ns_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m68_0_ns_1_LC_8_14_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.bcd2segment1.m68_0_ns_1_LC_8_14_1  (
            .in0(N__16883),
            .in1(N__13761),
            .in2(_gnd_net_),
            .in3(N__18902),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m68_0_ns_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m68_0_ns_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m68_0_ns_LC_8_14_2 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \Lab_UT.bcd2segment1.m68_0_ns_LC_8_14_2  (
            .in0(N__18960),
            .in1(N__13543),
            .in2(N__13596),
            .in3(N__13517),
            .lcout(\Lab_UT.m68_0_ns ),
            .ltout(\Lab_UT.m68_0_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIO00A3_3_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIO00A3_3_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIO00A3_3_LC_8_14_3 .LUT_INIT=16'b1111001011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIO00A3_3_LC_8_14_3  (
            .in0(N__13544),
            .in1(N__13593),
            .in2(N__13569),
            .in3(N__13566),
            .lcout(\Lab_UT.dictrl.next_state_set_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIFOTF_3_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIFOTF_3_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIFOTF_3_LC_8_14_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIFOTF_3_LC_8_14_4  (
            .in0(N__18901),
            .in1(N__18959),
            .in2(_gnd_net_),
            .in3(N__13542),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIB7JE1_1_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIB7JE1_1_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIB7JE1_1_LC_8_14_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIB7JE1_1_LC_8_14_5  (
            .in0(N__13518),
            .in1(_gnd_net_),
            .in2(N__13482),
            .in3(N__13731),
            .lcout(\Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_LC_8_14_6 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_2_LC_8_14_6  (
            .in0(N__17887),
            .in1(N__17307),
            .in2(N__13479),
            .in3(N__17520),
            .lcout(\Lab_UT.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18429),
            .ce(),
            .sr(N__18695));
    defparam \Lab_UT.dictrl.state_0_RNIEI8U_2_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIEI8U_2_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIEI8U_2_LC_8_14_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIEI8U_2_LC_8_14_7  (
            .in0(N__16882),
            .in1(N__13762),
            .in2(N__18967),
            .in3(N__18900),
            .lcout(\Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_3_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_3_0 .LUT_INIT=16'b1111100111100010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_3_0  (
            .in0(N__19350),
            .in1(N__19286),
            .in2(N__19182),
            .in3(N__19074),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_314_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_9_3_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_314_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13725),
            .in3(N__14976),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__18668));
    defparam \uu2.bitmap_87_LC_9_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_9_3_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_87_LC_9_3_4  (
            .in0(N__14978),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13722),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__18668));
    defparam \uu2.bitmap_RNI672H_84_LC_9_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI672H_84_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI672H_84_LC_9_3_5 .LUT_INIT=16'b0001010110011101;
    LogicCell40 \uu2.bitmap_RNI672H_84_LC_9_3_5  (
            .in0(N__13981),
            .in1(N__15050),
            .in2(N__13695),
            .in3(N__13707),
            .lcout(\uu2.m76_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_84_LC_9_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_9_3_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_84_LC_9_3_6  (
            .in0(N__14977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17589),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__18668));
    defparam \uu2.w_addr_displaying_fast_7_LC_9_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_9_3_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_9_3_7  (
            .in0(N__15310),
            .in1(N__15477),
            .in2(N__15397),
            .in3(N__15051),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__18668));
    defparam \uu2.bitmap_168_LC_9_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_9_4_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_168_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__13686),
            .in2(_gnd_net_),
            .in3(N__14986),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__18667));
    defparam \Lab_UT.bcd2segment1.m109_LC_9_4_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m109_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m109_LC_9_4_2 .LUT_INIT=16'b1110110011110010;
    LogicCell40 \Lab_UT.bcd2segment1.m109_LC_9_4_2  (
            .in0(N__14267),
            .in1(N__14178),
            .in2(N__14100),
            .in3(N__16262),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_72_LC_9_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_9_4_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_72_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13653),
            .in3(N__14988),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__18667));
    defparam \Lab_UT.bcd2segment1.m113_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m113_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m113_LC_9_4_4 .LUT_INIT=16'b1110111111101010;
    LogicCell40 \Lab_UT.bcd2segment1.m113_LC_9_4_4  (
            .in0(N__14268),
            .in1(N__14179),
            .in2(N__14101),
            .in3(N__16263),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.N_248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_200_LC_9_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_9_4_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_200_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14010),
            .in3(N__14987),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__18667));
    defparam \uu2.bitmap_RNI65TM_72_LC_9_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI65TM_72_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI65TM_72_LC_9_4_6 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \uu2.bitmap_RNI65TM_72_LC_9_4_6  (
            .in0(N__14007),
            .in1(N__15043),
            .in2(N__13985),
            .in3(N__14001),
            .lcout(\uu2.m76_bm_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_0_LC_9_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(N__13980),
            .in2(_gnd_net_),
            .in3(N__15470),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__18667));
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_9_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_9_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_26_LC_9_5_0  (
            .in0(N__15542),
            .in1(N__14621),
            .in2(N__15312),
            .in3(N__15112),
            .lcout(\uu2.mem0.g1_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_9_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_9_5_1 .LUT_INIT=16'b0101111001011010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_43_LC_9_5_1  (
            .in0(N__15113),
            .in1(N__15281),
            .in2(N__14650),
            .in3(N__15543),
            .lcout(\uu2.mem0.g2_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_9_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_9_5_2 .LUT_INIT=16'b0011001111101100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_63_LC_9_5_2  (
            .in0(N__15541),
            .in1(N__14620),
            .in2(N__15311),
            .in3(N__15111),
            .lcout(\uu2.mem0.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_9_5_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_9_5_3 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_68_LC_9_5_3  (
            .in0(N__13908),
            .in1(N__16119),
            .in2(_gnd_net_),
            .in3(N__13833),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_9_5_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_9_5_4 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_45_LC_9_5_4  (
            .in0(N__14731),
            .in1(_gnd_net_),
            .in2(N__14700),
            .in3(N__14691),
            .lcout(\uu2.mem0.bitmap_pmux_u_i_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_9_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_9_5_5 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_69_LC_9_5_5  (
            .in0(N__15110),
            .in1(N__15274),
            .in2(N__14649),
            .in3(N__15540),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_6_LC_9_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_9_5_6 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_9_5_6 .LUT_INIT=16'b1101010110101010;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_9_5_6  (
            .in0(N__15283),
            .in1(N__14625),
            .in2(N__15196),
            .in3(N__15374),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_ness_6C_net ),
            .ce(N__14580),
            .sr(N__18665));
    defparam \uu2.w_addr_displaying_nesr_8_LC_9_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_8_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_8_LC_9_5_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_nesr_8_LC_9_5_7  (
            .in0(N__15373),
            .in1(N__15179),
            .in2(N__14651),
            .in3(N__15282),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_ness_6C_net ),
            .ce(N__14580),
            .sr(N__18665));
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_49_LC_9_6_0  (
            .in0(N__14802),
            .in1(N__15309),
            .in2(N__15993),
            .in3(N__15538),
            .lcout(),
            .ltout(\uu2.mem0.G_13_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_6_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_6_1 .LUT_INIT=16'b0111000001000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_27_LC_9_6_1  (
            .in0(N__15672),
            .in1(N__15714),
            .in2(N__14544),
            .in3(N__14541),
            .lcout(),
            .ltout(\uu2.mem0.G_13_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_6_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_6_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_9_6_2  (
            .in0(N__14530),
            .in1(N__14421),
            .in2(N__14400),
            .in3(N__14384),
            .lcout(\uu2.mem0.G_13_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_86_LC_9_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_86_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_86_LC_9_6_3 .LUT_INIT=16'b0011001100000101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_86_LC_9_6_3  (
            .in0(N__15537),
            .in1(N__15977),
            .in2(N__14805),
            .in3(N__15259),
            .lcout(\uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI59BR1_5_LC_9_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI59BR1_5_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI59BR1_5_LC_9_6_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI59BR1_5_LC_9_6_4  (
            .in0(N__15715),
            .in1(N__15673),
            .in2(_gnd_net_),
            .in3(N__15539),
            .lcout(\uu2.N_12_i ),
            .ltout(\uu2.N_12_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_LC_9_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_rep1_LC_9_6_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_LC_9_6_5  (
            .in0(N__15476),
            .in1(N__15261),
            .in2(N__15720),
            .in3(N__15981),
            .lcout(\uu2.w_addr_displaying_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7_rep1C_net ),
            .ce(),
            .sr(N__18662));
    defparam \uu2.w_addr_displaying_5_LC_9_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_9_6_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_9_6_6  (
            .in0(N__15716),
            .in1(N__15674),
            .in2(N__15579),
            .in3(N__15474),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7_rep1C_net ),
            .ce(),
            .sr(N__18662));
    defparam \uu2.w_addr_displaying_7_LC_9_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_9_6_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_7_LC_9_6_7  (
            .in0(N__15475),
            .in1(N__15149),
            .in2(N__15386),
            .in3(N__15260),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7_rep1C_net ),
            .ce(),
            .sr(N__18662));
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_7_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNIKGSI_58_LC_9_7_1  (
            .in0(N__14997),
            .in1(N__15052),
            .in2(_gnd_net_),
            .in3(N__14823),
            .lcout(\uu2.N_272 ),
            .ltout(\uu2.N_272_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_9_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_9_7_2 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_52_LC_9_7_2  (
            .in0(N__14817),
            .in1(N__14804),
            .in2(N__15012),
            .in3(N__15009),
            .lcout(\uu2.mem0.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_58_LC_9_7_3 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_9_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_58_LC_9_7_3  (
            .in0(N__17607),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14975),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_58C_net ),
            .ce(),
            .sr(N__18661));
    defparam \uu2.bitmap_186_LC_9_7_5 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_9_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_186_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__17598),
            .in2(_gnd_net_),
            .in3(N__14974),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_58C_net ),
            .ce(),
            .sr(N__18661));
    defparam \uu2.mem0.ram512X8_inst_RNO_81_LC_9_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_81_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_81_LC_9_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_81_LC_9_7_6  (
            .in0(N__14816),
            .in1(N__14803),
            .in2(_gnd_net_),
            .in3(N__14742),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_9_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_9_7_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_56_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__16118),
            .in2(N__16050),
            .in3(N__16020),
            .lcout(\uu2.mem0.N_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_0_LC_9_8_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_0_LC_9_8_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_0_LC_9_8_0 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \buart.Z_rx.bitcount_0_LC_9_8_0  (
            .in0(N__17227),
            .in1(N__16563),
            .in2(N__17039),
            .in3(N__16511),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \buart.Z_rx.bitcount_4_LC_9_8_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_4_LC_9_8_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_4_LC_9_8_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \buart.Z_rx.bitcount_4_LC_9_8_1  (
            .in0(N__16510),
            .in1(N__17038),
            .in2(N__17273),
            .in3(N__16128),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \buart.Z_rx.bitcount_1_LC_9_8_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_1_LC_9_8_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_1_LC_9_8_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \buart.Z_rx.bitcount_1_LC_9_8_2  (
            .in0(N__16524),
            .in1(N__17449),
            .in2(N__17040),
            .in3(N__16512),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \buart.Z_rx.bitcount_2_LC_9_8_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_2_LC_9_8_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_2_LC_9_8_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \buart.Z_rx.bitcount_2_LC_9_8_3  (
            .in0(N__16509),
            .in1(N__17037),
            .in2(N__17182),
            .in3(N__16419),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \uu2.mem0.ram512X8_inst_RNO_80_LC_9_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_80_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_80_LC_9_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_80_LC_9_8_4  (
            .in0(N__15982),
            .in1(N__16037),
            .in2(_gnd_net_),
            .in3(N__16026),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_82_LC_9_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_82_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_82_LC_9_8_5 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_82_LC_9_8_5  (
            .in0(N__16007),
            .in1(N__15983),
            .in2(_gnd_net_),
            .in3(N__15917),
            .lcout(\uu2.mem0.N_98_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_2_LC_9_8_6 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_9_8_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_2_LC_9_8_6  (
            .in0(N__15795),
            .in1(N__15868),
            .in2(N__15849),
            .in3(N__15737),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \uu2.r_addr_1_LC_9_8_7 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_9_8_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_1_LC_9_8_7  (
            .in0(N__15736),
            .in1(N__15844),
            .in2(_gnd_net_),
            .in3(N__15794),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18476),
            .ce(),
            .sr(N__18692));
    defparam \Lab_UT.didp.ce_1_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_9_9_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_9_9_0  (
            .in0(N__19069),
            .in1(N__19367),
            .in2(N__19177),
            .in3(N__19281),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18468),
            .ce(),
            .sr(N__18235));
    defparam \Lab_UT.bcd2segment1.m53_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m53_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m53_LC_9_9_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Lab_UT.bcd2segment1.m53_LC_9_9_1  (
            .in0(N__16832),
            .in1(N__19068),
            .in2(_gnd_net_),
            .in3(N__16397),
            .lcout(\Lab_UT.bcd2segment1.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_2_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_9_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_9_9_3  (
            .in0(N__18822),
            .in1(N__19434),
            .in2(N__18111),
            .in3(N__18095),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18468),
            .ce(),
            .sr(N__18235));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__16279),
            .in2(_gnd_net_),
            .in3(N__16253),
            .lcout(\Lab_UT.didp.countrce3.q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_10_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__17230),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_10_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__17453),
            .in2(_gnd_net_),
            .in3(N__16155),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_10_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17197),
            .in3(N__16152),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_10_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17415),
            .in3(N__16134),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_10_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_4_LC_9_10_4  (
            .in0(N__17366),
            .in1(N__16491),
            .in2(N__17274),
            .in3(N__16131),
            .lcout(\buart.Z_rx.bitcount_lm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m42_bm_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m42_bm_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m42_bm_LC_9_10_6 .LUT_INIT=16'b0011101100001011;
    LogicCell40 \Lab_UT.bcd2segment1.m42_bm_LC_9_10_6  (
            .in0(N__16848),
            .in1(N__16821),
            .in2(N__16728),
            .in3(N__18180),
            .lcout(\Lab_UT.bcd2segment1.m42_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_9_10_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_9_10_7 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_0_LC_9_10_7  (
            .in0(N__16490),
            .in1(N__16599),
            .in2(N__17235),
            .in3(N__17367),
            .lcout(\buart.Z_rx.bitcount_lm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_RNIMK771_4_LC_9_11_0  (
            .in0(N__17451),
            .in1(N__17269),
            .in2(N__17198),
            .in3(N__17409),
            .lcout(),
            .ltout(\buart.Z_rx.un1_sample_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_9_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_9_11_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIC77M1_0_LC_9_11_1  (
            .in0(N__17098),
            .in1(N__17127),
            .in2(N__16554),
            .in3(N__17234),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_9_11_2 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_3_LC_9_11_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_9_11_2  (
            .in0(N__16972),
            .in1(N__17006),
            .in2(N__17561),
            .in3(N__16938),
            .lcout(\Lab_UT.dictrl.next_state_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18454),
            .ce(N__17495),
            .sr(N__16542));
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_9_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_9_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIAPJJ_1_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__17404),
            .in2(_gnd_net_),
            .in3(N__17450),
            .lcout(\buart.Z_rx.idle_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_11_6 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_1_LC_9_11_6  (
            .in0(N__17452),
            .in1(N__16530),
            .in2(N__17373),
            .in3(N__16488),
            .lcout(\buart.Z_rx.bitcount_lm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_11_7 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_2_LC_9_11_7  (
            .in0(N__16489),
            .in1(N__16425),
            .in2(N__17199),
            .in3(N__17372),
            .lcout(\buart.Z_rx.bitcount_lm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_2_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_9_12_0 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_2_LC_9_12_0 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_9_12_0  (
            .in0(N__17298),
            .in1(N__17338),
            .in2(N__17565),
            .in3(N__17529),
            .lcout(\Lab_UT.dictrl.next_state_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18447),
            .ce(N__17496),
            .sr(N__17472));
    defparam \buart.Z_rx.bitcount_RNIBQJJ_4_LC_9_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIBQJJ_4_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIBQJJ_4_LC_9_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIBQJJ_4_LC_9_12_1  (
            .in0(N__17454),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17268),
            .lcout(),
            .ltout(\buart.Z_rx.valid_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_9_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_9_12_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_0_LC_9_12_2  (
            .in0(N__17186),
            .in1(N__17229),
            .in2(N__17418),
            .in3(N__17405),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_9_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_9_12_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \buart.Z_rx.bitcount_RNIIU223_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17376),
            .in3(N__17138),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI9T1T1_2_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI9T1T1_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI9T1T1_2_LC_9_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI9T1T1_2_LC_9_12_5  (
            .in0(N__17337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17313),
            .lcout(\Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_9_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_9_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_4_LC_9_12_6  (
            .in0(N__17267),
            .in1(N__17228),
            .in2(N__17196),
            .in3(N__17145),
            .lcout(\buart.Z_rx.idle ),
            .ltout(\buart.Z_rx.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_9_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_9_12_7 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \buart.Z_rx.bitcount_RNILM873_0_LC_9_12_7  (
            .in0(N__17123),
            .in1(N__17099),
            .in2(N__17061),
            .in3(N__17054),
            .lcout(\buart.Z_rx.bitcountlde_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_LC_9_13_4 .LUT_INIT=16'b1010001111110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_LC_9_13_4  (
            .in0(N__17010),
            .in1(N__16976),
            .in2(N__17895),
            .in3(N__16935),
            .lcout(\Lab_UT.state_i_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18440),
            .ce(),
            .sr(N__18696));
    defparam \Lab_UT.dictrl.state_ret_1_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_LC_9_13_6 .LUT_INIT=16'b1010001111110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_LC_9_13_6  (
            .in0(N__17947),
            .in1(N__17919),
            .in2(N__17894),
            .in3(N__17805),
            .lcout(\Lab_UT.state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18440),
            .ce(),
            .sr(N__18696));
    defparam \buart.Z_rx.shifter_2_LC_9_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17756),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18434),
            .ce(N__17652),
            .sr(N__18713));
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_11_7_0 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_0_LC_11_7_0  (
            .in0(N__19313),
            .in1(N__19226),
            .in2(N__19141),
            .in3(N__19024),
            .lcout(\Lab_UT.bcd2segment1.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m96_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m96_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m96_LC_11_7_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \Lab_UT.bcd2segment1.m96_LC_11_7_4  (
            .in0(N__19312),
            .in1(N__19227),
            .in2(N__19140),
            .in3(N__19025),
            .lcout(\Lab_UT.bcd2segment1.N_192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_11_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_11_8_0  (
            .in0(N__18796),
            .in1(N__18844),
            .in2(_gnd_net_),
            .in3(N__19038),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_11_8_1 .LUT_INIT=16'b1111101111000010;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_5_LC_11_8_1  (
            .in0(N__18080),
            .in1(N__19422),
            .in2(N__18017),
            .in3(N__18159),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_11_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_11_8_2 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_11_8_2  (
            .in0(N__18797),
            .in1(N__19039),
            .in2(N__19264),
            .in3(N__18845),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_11_8_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_11_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.bcd2segment2.un1_num_5_2_LC_11_8_3  (
            .in0(N__18083),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18160),
            .lcout(\Lab_UT.three_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_11_8_4 .LUT_INIT=16'b1111100111100010;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_3_LC_11_8_4  (
            .in0(N__19424),
            .in1(N__18157),
            .in2(N__18019),
            .in3(N__18082),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_11_8_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_11_8_5 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_4_LC_11_8_5  (
            .in0(N__18081),
            .in1(N__19423),
            .in2(N__18018),
            .in3(N__18158),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m1_LC_11_8_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m1_LC_11_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m1_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__19243),
            .in2(_gnd_net_),
            .in3(N__19037),
            .lcout(),
            .ltout(\Lab_UT.three_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_11_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_11_8_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_11_8_7  (
            .in0(N__18846),
            .in1(N__18798),
            .in2(N__18183),
            .in3(N__19329),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_9_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_11_9_0  (
            .in0(N__18085),
            .in1(N__18522),
            .in2(_gnd_net_),
            .in3(N__19467),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18478),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_11_9_1 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_11_9_1  (
            .in0(N__18162),
            .in1(N__18526),
            .in2(N__19473),
            .in3(N__18086),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18478),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI4V78_3_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI4V78_3_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI4V78_3_LC_11_9_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI4V78_3_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__18015),
            .in2(_gnd_net_),
            .in3(N__18161),
            .lcout(\Lab_UT.didp.countrce2.un15_ce_2 ),
            .ltout(\Lab_UT.didp.countrce2.un15_ce_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_2_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_2_LC_11_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI84NN1_2_LC_11_9_3  (
            .in0(N__18814),
            .in1(N__19428),
            .in2(N__18099),
            .in3(N__18084),
            .lcout(\Lab_UT.q_RNI84NN1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_11_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__19451),
            .in2(_gnd_net_),
            .in3(N__19429),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_11_9_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_11_9_6  (
            .in0(N__18527),
            .in1(N__19468),
            .in2(N__18030),
            .in3(N__18016),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18478),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_11_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_11_9_7 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_11_9_7  (
            .in0(N__19472),
            .in1(N__19452),
            .in2(N__18528),
            .in3(N__19430),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18478),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_11_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_11_10_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_11_10_1  (
            .in0(N__19054),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__19260),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_11_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_11_10_2 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_11_10_2  (
            .in0(N__19115),
            .in1(N__18795),
            .in2(N__19371),
            .in3(N__18843),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18470),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.m5_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.m5_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.m5_LC_11_10_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.bcd2segment1.m5_LC_11_10_6  (
            .in0(N__19338),
            .in1(N__19256),
            .in2(N__19136),
            .in3(N__19053),
            .lcout(\Lab_UT.nine ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_0_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_11_11_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_11_11_0  (
            .in0(N__18987),
            .in1(N__18968),
            .in2(_gnd_net_),
            .in3(N__18909),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18461),
            .ce(),
            .sr(N__18246));
    defparam \Lab_UT.didp.reset_0_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_0_LC_11_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.reset_0_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__18815),
            .in2(_gnd_net_),
            .in3(N__18750),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18461),
            .ce(),
            .sr(N__18246));
    defparam \Lab_UT.didp.reset_1_LC_12_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_1_LC_12_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.reset_1_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__18766),
            .in2(_gnd_net_),
            .in3(N__18749),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18486),
            .ce(),
            .sr(N__18242));
endmodule // latticehx1k
