-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 21 2019 00:12:19

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__22472\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.un143_ci_0_cascade_\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.un4_l_count_16_cascade_\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \buart.Z_rx.idle_0_cascade_\ : std_logic;
signal \buart.Z_rx.valid_0_cascade_\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \buart.Z_rx.N_27_0_i_cascade_\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3_cascade_\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un165_ci_0_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un187_ci_1\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un44_ci\ : std_logic;
signal \uu0.un44_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \resetGen.reset_count_2_0_4\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.un404_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.N_34\ : std_logic;
signal \uu2.N_34_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.N_31\ : std_logic;
signal \uu2.N_31_cascade_\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.didp.regrce3.LdAMones_0\ : std_logic;
signal \G_184\ : std_logic;
signal \G_184_cascade_\ : std_logic;
signal \Lab_UT.un1_idle_1_0_iclkZ0_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_117_cascade_\ : std_logic;
signal \G_180_cascade_\ : std_logic;
signal \G_181_cascade_\ : std_logic;
signal \G_180\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_0_cascade_\ : std_logic;
signal \G_179_cascade_\ : std_logic;
signal \Lab_UT.alarmstate_0_sqmuxa_1\ : std_logic;
signal \Lab_UT.un1_idle_5_0_iclkZ0_cascade_\ : std_logic;
signal \Lab_UT.un1_armed_2_0_iso_iZ0\ : std_logic;
signal \G_185\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu2.un28_w_addr_user_i_cascade_\ : std_logic;
signal \uu2.un51_w_data_displaying_i_a2_1\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a3_2_0\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_3C_net\ : std_logic;
signal \uu2.w_addr_displaying_RNI03P31Z0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \uu2.N_406_cascade_\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \uu2.N_383_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\ : std_logic;
signal \uu2.bitmap_pmux_u_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\ : std_logic;
signal \uu2.w_addr_displaying_RNI0NG56Z0Z_4\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4_cascade_\ : std_logic;
signal \uu2.un20_w_addr_userZ0Z_1\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_3\ : std_logic;
signal \Lab_UT.dispString.N_140\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \G_188\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_3\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \G_186_cascade_\ : std_logic;
signal \G_187\ : std_logic;
signal \G_187_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_1_iv_i_1_4\ : std_logic;
signal \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \G_182\ : std_logic;
signal \G_183\ : std_logic;
signal \G_182_cascade_\ : std_logic;
signal \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z8\ : std_logic;
signal \Lab_UT.dictrl.g1_0_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_5_4_0_cascade_\ : std_logic;
signal \uu2.un28_w_addr_user_i\ : std_logic;
signal \INVuu2.w_addr_user_2C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i5_mux\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15_cascade_\ : std_logic;
signal \uu2.N_401\ : std_logic;
signal \INVuu2.w_addr_displaying_1_rep1_nesrC_net\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \INVuu2.bitmap_197C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \Lab_UT.didp.ce_12_1\ : std_logic;
signal \Lab_UT.didp.ce_12_1_cascade_\ : std_logic;
signal \Lab_UT.didp.ce_12_3_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.ce_12_1_1\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3\ : std_logic;
signal \Lab_UT.dispString.N_137\ : std_logic;
signal \uu0_sec_clkD\ : std_logic;
signal \Lab_UT.dispString.N_143_cascade_\ : std_logic;
signal \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.dispString.un42_dOutP_1\ : std_logic;
signal \Lab_UT.dispString.N_102_cascade_\ : std_logic;
signal \G_186\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_4\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_3\ : std_logic;
signal \G_179\ : std_logic;
signal \G_181\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_144\ : std_logic;
signal \Lab_UT.dispString.N_124\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_95\ : std_logic;
signal \Lab_UT.dispString.N_102\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \Lab_UT.dispString.N_143\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_1_1\ : std_logic;
signal \Lab_UT.didp.regrce2.LdAStens_0\ : std_logic;
signal \Lab_UT.dictrl.g1_4_0\ : std_logic;
signal \Lab_UT.dictrl.g1_5_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_5_3_0\ : std_logic;
signal \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\ : std_logic;
signal \resetGen.escKeyZ0Z_4_cascade_\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \resetGen.escKeyZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.g1_0Z0Z_5\ : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_8C_net\ : std_logic;
signal \uu2.N_37\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_36\ : std_logic;
signal \INVuu2.bitmap_40C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \uu2.N_14_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux\ : std_logic;
signal \uu2.bitmap_RNI2Q8F1Z0Z_111\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.N_24_cascade_\ : std_logic;
signal \uu2.N_31_i\ : std_logic;
signal \uu2.N_166\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1_cascade_\ : std_logic;
signal \uu2.N_26\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.N_149\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.N_25\ : std_logic;
signal \Lab_UT.didp.un24_ce_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.N_96\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.didp.regrce4.LdAMtens_0\ : std_logic;
signal \Lab_UT.dispString.N_145\ : std_logic;
signal \Lab_UT.dispString.N_118_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_i_0_1\ : std_logic;
signal \Lab_UT.didp.regrce1.LdASones_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_4\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_o3_5\ : std_logic;
signal \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_11_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_0\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_a5_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_18_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_6_3_0\ : std_logic;
signal \Lab_UT.dictrl.g2Z0Z_0\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.dictrl.g1_1_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_1_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.N_3\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m37_N_2LZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux_1\ : std_logic;
signal \Lab_UT.i8_mux_0_cascade_\ : std_logic;
signal \Lab_UT.didp.g0_0_2Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_sn\ : std_logic;
signal \Lab_UT.dictrl.g1_1_0_1_cascade_\ : std_logic;
signal \Lab_UT.g1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_rn_0\ : std_logic;
signal \Lab_UT.dictrl.m22Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_3_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux_0\ : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal \uu2.N_40\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.N_45\ : std_logic;
signal \INVuu2.w_addr_displaying_ness_6C_net\ : std_logic;
signal \uu2.N_33_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \INVuu2.w_addr_displaying_7C_net\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.didp.reset_12_1_3\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.didp.countrce2.N_93\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.sec1_1\ : std_logic;
signal \Lab_UT.sec1_2\ : std_logic;
signal \Lab_UT.sec1_3\ : std_logic;
signal \Lab_UT.sec1_0\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \uu2.bitmap_pmux_17_ns_1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.bitmap_pmux_16_ns_1\ : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_8\ : std_logic;
signal \uu2.N_44\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \Lab_UT.min2_2\ : std_logic;
signal \Lab_UT.min2_3\ : std_logic;
signal \Lab_UT.min2_0\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \INVuu2.bitmap_215C_net\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.min2_1\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMtens_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMones_1\ : std_logic;
signal \Lab_UT.LdAMones\ : std_logic;
signal \Lab_UT.LdAMones_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_2_fast\ : std_logic;
signal \Lab_UT.dictrl.dicRun_1\ : std_logic;
signal \Lab_UT.LdASones\ : std_logic;
signal \Lab_UT.LdAStens\ : std_logic;
signal \Lab_UT.dictrl.N_22\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_20_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_22_0_0\ : std_logic;
signal \Lab_UT.didp.g0_0Z0Z_2\ : std_logic;
signal \Lab_UT.next_state_1_0_0_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state6\ : std_logic;
signal \Lab_UT.dictrl.m19_1\ : std_logic;
signal \Lab_UT.dictrl.m19_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_20\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_20_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_4_2\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_0\ : std_logic;
signal \Lab_UT.dictrl.g2_0_0\ : std_logic;
signal \shifter_1_rep1_RNI0FPF\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_1\ : std_logic;
signal \N_15\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_1_cascade_\ : std_logic;
signal \N_14_0\ : std_logic;
signal \Lab_UT.dictrl.N_20_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state66_2\ : std_logic;
signal \Lab_UT.dictrl.state_i_3_0\ : std_logic;
signal \N_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_67_mux\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_12\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g0_3_4\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m22_xZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_72_mux_cascade_\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal \Lab_UT.dictrl.m34Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g1_0_xZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0_4\ : std_logic;
signal \Lab_UT.dictrl.g0_5_3\ : std_logic;
signal \Lab_UT.dictrl.g1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m22Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.g0_5Z0Z_4\ : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal \G_6_0_a6_3_3\ : std_logic;
signal \buart__rx_shifter_fast_4\ : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.un3_w_addr_user_4_cascade_\ : std_logic;
signal \uu2.un3_w_addr_user_5\ : std_logic;
signal \uu2.un3_w_addr_user\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.un426_ci_3\ : std_logic;
signal \uu2.un404_ci_cascade_\ : std_logic;
signal \uu2.vbuf_w_addr_user.un448_ci_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.w_addr_user_RNI43E87Z0Z_4\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmap_pmux_20_ns_1\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.bitmap_pmux_26_bm_1\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.bitmap_RNIP2JO1Z0Z_34\ : std_logic;
signal \Lab_UT.min1_0\ : std_logic;
signal \Lab_UT.min1_3\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmap_pmux_19_ns_1\ : std_logic;
signal \Lab_UT.sec2_0\ : std_logic;
signal \Lab_UT.sec2_3\ : std_logic;
signal \Lab_UT.sec2_1\ : std_logic;
signal \Lab_UT.sec2_2\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \uu2.bitmap_RNIM5E21Z0Z_314\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \uu2.N_152\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.min1_1\ : std_logic;
signal \Lab_UT.didp.countrce4.un13_qPone\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3\ : std_logic;
signal \Lab_UT.didp.countrce1.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.loadalarm_0\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.min1_2\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.state_ret_8_ess\ : std_logic;
signal \Lab_UT.next_state_0\ : std_logic;
signal \Lab_UT.didp.N_90\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.LdSones_i_4\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_rn_0\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_57_1\ : std_logic;
signal \Lab_UT.dictrl.N_55_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_2\ : std_logic;
signal \Lab_UT.bu_rx_data_rdy_0\ : std_logic;
signal \Lab_UT.dictrl.g0_1_mb_sn\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_1\ : std_logic;
signal \Lab_UT.dictrl.un15_loadalarm_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.loadalarm_0_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \Lab_UT.next_state_1\ : std_logic;
signal \Lab_UT.next_state_2\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.dictrl.m34_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.N_33_0\ : std_logic;
signal \Lab_UT.dictrl.N_60_0_0\ : std_logic;
signal \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_26_0\ : std_logic;
signal \Lab_UT.dictrl.i8_mux_0\ : std_logic;
signal \Lab_UT.dictrl.m34_0\ : std_logic;
signal \Lab_UT.dictrl.N_18\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_3\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.g0_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0\ : std_logic;
signal \Lab_UT.un1_next_state66_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\ : std_logic;
signal m7_a0 : std_logic;
signal \Lab_UT.dictrl.N_8_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_0_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_6_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_8_0\ : std_logic;
signal \Lab_UT.dictrl.i9_mux\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.N_60\ : std_logic;
signal \Lab_UT.dictrl.i8_mux_cascade_\ : std_logic;
signal \Lab_UT.dicLdSones_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_0Z0Z_0\ : std_logic;
signal \Lab_UT.stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_59\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal \Lab_UT.dictrl.N_15_0\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_3_rep2 : std_logic;
signal \G_6_0_a6_2\ : std_logic;
signal \Lab_UT.dictrl.state_0_rep1\ : std_logic;
signal \N_63_mux\ : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \Lab_UT.dictrl.N_72_mux\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m13_out\ : std_logic;
signal \Lab_UT.dictrl.N_59_1_0\ : std_logic;
signal \Lab_UT.dictrl.state_fast_0\ : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \Lab_UT.dictrl.g1_1Z0Z_5\ : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal \Lab_UT.dictrl.g1_1_4_cascade_\ : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0\ : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal \Lab_UT.dictrl.g0_6_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_57_0\ : std_logic;
signal \Lab_UT.dictrl.g0_6_3\ : std_logic;
signal \Lab_UT.dictrl.g1_1\ : std_logic;
signal \Lab_UT.dictrl.gZ0Z2\ : std_logic;
signal \Lab_UT_dictrl_state_1\ : std_logic;
signal \Lab_UT.dictrl.N_55_0\ : std_logic;
signal \Lab_UT.state_i_4_3\ : std_logic;
signal \Lab_UT.dictrl.g1_rn_0_cascade_\ : std_logic;
signal \Lab_UT.state_2\ : std_logic;
signal \Lab_UT.dictrl.G_25_i_a5_1_0_0\ : std_logic;
signal rst_g : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c2\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal clk_g : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__9865\&\N__9850\&\N__9805\&\N__10116\&\N__10207\&\N__9832\&\N__9928\&\N__9901\&\N__10261\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__10417\&\N__13063\&\N__13192\&\N__13075\&\N__13123\&\N__16063\&\N__21733\&\N__20644\&\N__9247\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__9775\&'0'&\N__9979\&'0'&\N__9952\&'0'&\N__9964\&'0'&\N__10219\&'0'&\N__9958\&'0'&\N__9934\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__8074\,
            RESETB => \N__10849\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22345\,
            RE => \N__10845\,
            WCLKE => \N__10608\,
            WCLK => \N__22344\,
            WE => \N__10609\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22472\,
            DIN => \N__22471\,
            DOUT => \N__22470\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22472\,
            PADOUT => \N__22471\,
            PADIN => \N__22470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22463\,
            DIN => \N__22462\,
            DOUT => \N__22461\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22463\,
            PADOUT => \N__22462\,
            PADIN => \N__22461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22454\,
            DIN => \N__22453\,
            DOUT => \N__22452\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22454\,
            PADOUT => \N__22453\,
            PADIN => \N__22452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22445\,
            DIN => \N__22444\,
            DOUT => \N__22443\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__22445\,
            PADOUT => \N__22444\,
            PADIN => \N__22443\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__22299\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22436\,
            DIN => \N__22435\,
            DOUT => \N__22434\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22436\,
            PADOUT => \N__22435\,
            PADIN => \N__22434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22427\,
            DIN => \N__22426\,
            DOUT => \N__22425\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22427\,
            PADOUT => \N__22426\,
            PADIN => \N__22425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22418\,
            DIN => \N__22417\,
            DOUT => \N__22416\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22418\,
            PADOUT => \N__22417\,
            PADIN => \N__22416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22409\,
            DIN => \N__22408\,
            DOUT => \N__22407\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22409\,
            PADOUT => \N__22408\,
            PADIN => \N__22407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22400\,
            DIN => \N__22399\,
            DOUT => \N__22398\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22400\,
            PADOUT => \N__22399\,
            PADIN => \N__22398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8392\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22391\,
            DIN => \N__22390\,
            DOUT => \N__22389\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22391\,
            PADOUT => \N__22390\,
            PADIN => \N__22389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5450\ : InMux
    port map (
            O => \N__22372\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__5449\ : InMux
    port map (
            O => \N__22369\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__5448\ : InMux
    port map (
            O => \N__22366\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__5447\ : InMux
    port map (
            O => \N__22363\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__5446\ : InMux
    port map (
            O => \N__22360\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__5444\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__22351\,
            I => \N__22260\
        );

    \I__5442\ : ClkMux
    port map (
            O => \N__22350\,
            I => \N__22081\
        );

    \I__5441\ : ClkMux
    port map (
            O => \N__22349\,
            I => \N__22081\
        );

    \I__5440\ : ClkMux
    port map (
            O => \N__22348\,
            I => \N__22081\
        );

    \I__5439\ : ClkMux
    port map (
            O => \N__22347\,
            I => \N__22081\
        );

    \I__5438\ : ClkMux
    port map (
            O => \N__22346\,
            I => \N__22081\
        );

    \I__5437\ : ClkMux
    port map (
            O => \N__22345\,
            I => \N__22081\
        );

    \I__5436\ : ClkMux
    port map (
            O => \N__22344\,
            I => \N__22081\
        );

    \I__5435\ : ClkMux
    port map (
            O => \N__22343\,
            I => \N__22081\
        );

    \I__5434\ : ClkMux
    port map (
            O => \N__22342\,
            I => \N__22081\
        );

    \I__5433\ : ClkMux
    port map (
            O => \N__22341\,
            I => \N__22081\
        );

    \I__5432\ : ClkMux
    port map (
            O => \N__22340\,
            I => \N__22081\
        );

    \I__5431\ : ClkMux
    port map (
            O => \N__22339\,
            I => \N__22081\
        );

    \I__5430\ : ClkMux
    port map (
            O => \N__22338\,
            I => \N__22081\
        );

    \I__5429\ : ClkMux
    port map (
            O => \N__22337\,
            I => \N__22081\
        );

    \I__5428\ : ClkMux
    port map (
            O => \N__22336\,
            I => \N__22081\
        );

    \I__5427\ : ClkMux
    port map (
            O => \N__22335\,
            I => \N__22081\
        );

    \I__5426\ : ClkMux
    port map (
            O => \N__22334\,
            I => \N__22081\
        );

    \I__5425\ : ClkMux
    port map (
            O => \N__22333\,
            I => \N__22081\
        );

    \I__5424\ : ClkMux
    port map (
            O => \N__22332\,
            I => \N__22081\
        );

    \I__5423\ : ClkMux
    port map (
            O => \N__22331\,
            I => \N__22081\
        );

    \I__5422\ : ClkMux
    port map (
            O => \N__22330\,
            I => \N__22081\
        );

    \I__5421\ : ClkMux
    port map (
            O => \N__22329\,
            I => \N__22081\
        );

    \I__5420\ : ClkMux
    port map (
            O => \N__22328\,
            I => \N__22081\
        );

    \I__5419\ : ClkMux
    port map (
            O => \N__22327\,
            I => \N__22081\
        );

    \I__5418\ : ClkMux
    port map (
            O => \N__22326\,
            I => \N__22081\
        );

    \I__5417\ : ClkMux
    port map (
            O => \N__22325\,
            I => \N__22081\
        );

    \I__5416\ : ClkMux
    port map (
            O => \N__22324\,
            I => \N__22081\
        );

    \I__5415\ : ClkMux
    port map (
            O => \N__22323\,
            I => \N__22081\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__22322\,
            I => \N__22081\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__22321\,
            I => \N__22081\
        );

    \I__5412\ : ClkMux
    port map (
            O => \N__22320\,
            I => \N__22081\
        );

    \I__5411\ : ClkMux
    port map (
            O => \N__22319\,
            I => \N__22081\
        );

    \I__5410\ : ClkMux
    port map (
            O => \N__22318\,
            I => \N__22081\
        );

    \I__5409\ : ClkMux
    port map (
            O => \N__22317\,
            I => \N__22081\
        );

    \I__5408\ : ClkMux
    port map (
            O => \N__22316\,
            I => \N__22081\
        );

    \I__5407\ : ClkMux
    port map (
            O => \N__22315\,
            I => \N__22081\
        );

    \I__5406\ : ClkMux
    port map (
            O => \N__22314\,
            I => \N__22081\
        );

    \I__5405\ : ClkMux
    port map (
            O => \N__22313\,
            I => \N__22081\
        );

    \I__5404\ : ClkMux
    port map (
            O => \N__22312\,
            I => \N__22081\
        );

    \I__5403\ : ClkMux
    port map (
            O => \N__22311\,
            I => \N__22081\
        );

    \I__5402\ : ClkMux
    port map (
            O => \N__22310\,
            I => \N__22081\
        );

    \I__5401\ : ClkMux
    port map (
            O => \N__22309\,
            I => \N__22081\
        );

    \I__5400\ : ClkMux
    port map (
            O => \N__22308\,
            I => \N__22081\
        );

    \I__5399\ : ClkMux
    port map (
            O => \N__22307\,
            I => \N__22081\
        );

    \I__5398\ : ClkMux
    port map (
            O => \N__22306\,
            I => \N__22081\
        );

    \I__5397\ : ClkMux
    port map (
            O => \N__22305\,
            I => \N__22081\
        );

    \I__5396\ : ClkMux
    port map (
            O => \N__22304\,
            I => \N__22081\
        );

    \I__5395\ : ClkMux
    port map (
            O => \N__22303\,
            I => \N__22081\
        );

    \I__5394\ : ClkMux
    port map (
            O => \N__22302\,
            I => \N__22081\
        );

    \I__5393\ : ClkMux
    port map (
            O => \N__22301\,
            I => \N__22081\
        );

    \I__5392\ : ClkMux
    port map (
            O => \N__22300\,
            I => \N__22081\
        );

    \I__5391\ : ClkMux
    port map (
            O => \N__22299\,
            I => \N__22081\
        );

    \I__5390\ : ClkMux
    port map (
            O => \N__22298\,
            I => \N__22081\
        );

    \I__5389\ : ClkMux
    port map (
            O => \N__22297\,
            I => \N__22081\
        );

    \I__5388\ : ClkMux
    port map (
            O => \N__22296\,
            I => \N__22081\
        );

    \I__5387\ : ClkMux
    port map (
            O => \N__22295\,
            I => \N__22081\
        );

    \I__5386\ : ClkMux
    port map (
            O => \N__22294\,
            I => \N__22081\
        );

    \I__5385\ : ClkMux
    port map (
            O => \N__22293\,
            I => \N__22081\
        );

    \I__5384\ : ClkMux
    port map (
            O => \N__22292\,
            I => \N__22081\
        );

    \I__5383\ : ClkMux
    port map (
            O => \N__22291\,
            I => \N__22081\
        );

    \I__5382\ : ClkMux
    port map (
            O => \N__22290\,
            I => \N__22081\
        );

    \I__5381\ : ClkMux
    port map (
            O => \N__22289\,
            I => \N__22081\
        );

    \I__5380\ : ClkMux
    port map (
            O => \N__22288\,
            I => \N__22081\
        );

    \I__5379\ : ClkMux
    port map (
            O => \N__22287\,
            I => \N__22081\
        );

    \I__5378\ : ClkMux
    port map (
            O => \N__22286\,
            I => \N__22081\
        );

    \I__5377\ : ClkMux
    port map (
            O => \N__22285\,
            I => \N__22081\
        );

    \I__5376\ : ClkMux
    port map (
            O => \N__22284\,
            I => \N__22081\
        );

    \I__5375\ : ClkMux
    port map (
            O => \N__22283\,
            I => \N__22081\
        );

    \I__5374\ : ClkMux
    port map (
            O => \N__22282\,
            I => \N__22081\
        );

    \I__5373\ : ClkMux
    port map (
            O => \N__22281\,
            I => \N__22081\
        );

    \I__5372\ : ClkMux
    port map (
            O => \N__22280\,
            I => \N__22081\
        );

    \I__5371\ : ClkMux
    port map (
            O => \N__22279\,
            I => \N__22081\
        );

    \I__5370\ : ClkMux
    port map (
            O => \N__22278\,
            I => \N__22081\
        );

    \I__5369\ : ClkMux
    port map (
            O => \N__22277\,
            I => \N__22081\
        );

    \I__5368\ : ClkMux
    port map (
            O => \N__22276\,
            I => \N__22081\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22275\,
            I => \N__22081\
        );

    \I__5366\ : ClkMux
    port map (
            O => \N__22274\,
            I => \N__22081\
        );

    \I__5365\ : ClkMux
    port map (
            O => \N__22273\,
            I => \N__22081\
        );

    \I__5364\ : ClkMux
    port map (
            O => \N__22272\,
            I => \N__22081\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22271\,
            I => \N__22081\
        );

    \I__5362\ : ClkMux
    port map (
            O => \N__22270\,
            I => \N__22081\
        );

    \I__5361\ : ClkMux
    port map (
            O => \N__22269\,
            I => \N__22081\
        );

    \I__5360\ : ClkMux
    port map (
            O => \N__22268\,
            I => \N__22081\
        );

    \I__5359\ : ClkMux
    port map (
            O => \N__22267\,
            I => \N__22081\
        );

    \I__5358\ : ClkMux
    port map (
            O => \N__22266\,
            I => \N__22081\
        );

    \I__5357\ : ClkMux
    port map (
            O => \N__22265\,
            I => \N__22081\
        );

    \I__5356\ : ClkMux
    port map (
            O => \N__22264\,
            I => \N__22081\
        );

    \I__5355\ : ClkMux
    port map (
            O => \N__22263\,
            I => \N__22081\
        );

    \I__5354\ : Glb2LocalMux
    port map (
            O => \N__22260\,
            I => \N__22081\
        );

    \I__5353\ : GlobalMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__5352\ : gio2CtrlBuf
    port map (
            O => \N__22078\,
            I => clk_g
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__5350\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22066\
        );

    \I__5349\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22066\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__22066\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__5346\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22054\
        );

    \I__5345\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22054\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22054\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__5343\ : CascadeMux
    port map (
            O => \N__22051\,
            I => \N__22047\
        );

    \I__5342\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22044\
        );

    \I__5341\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22041\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__22044\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__22041\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__5338\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22030\
        );

    \I__5337\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22030\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__22030\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__5335\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22022\
        );

    \I__5334\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22017\
        );

    \I__5333\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22017\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22022\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22017\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__22012\,
            I => \N__22007\
        );

    \I__5329\ : InMux
    port map (
            O => \N__22011\,
            I => \N__22001\
        );

    \I__5328\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22001\
        );

    \I__5327\ : InMux
    port map (
            O => \N__22007\,
            I => \N__21996\
        );

    \I__5326\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21996\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__22001\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__21996\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \N__21987\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__21990\,
            I => \N__21984\
        );

    \I__5321\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21979\
        );

    \I__5320\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21979\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__21979\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__5318\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21973\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__21973\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__5316\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21960\
        );

    \I__5315\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21960\
        );

    \I__5314\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21960\
        );

    \I__5313\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21957\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__21960\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__21957\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__21952\,
            I => \N__21948\
        );

    \I__5309\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21942\
        );

    \I__5308\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21935\
        );

    \I__5307\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21935\
        );

    \I__5306\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21935\
        );

    \I__5305\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21932\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__21942\,
            I => \N__21929\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21926\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__21932\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5301\ : Odrv12
    port map (
            O => \N__21929\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__21926\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__21919\,
            I => \N__21914\
        );

    \I__5298\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21904\
        );

    \I__5297\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21904\
        );

    \I__5296\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21886\
        );

    \I__5295\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21886\
        );

    \I__5294\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21886\
        );

    \I__5293\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21886\
        );

    \I__5292\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21886\
        );

    \I__5291\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21886\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21882\
        );

    \I__5289\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21879\
        );

    \I__5288\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21874\
        );

    \I__5287\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21874\
        );

    \I__5286\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21869\
        );

    \I__5285\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21869\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__21886\,
            I => \N__21863\
        );

    \I__5283\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21860\
        );

    \I__5282\ : Span4Mux_s2_h
    port map (
            O => \N__21882\,
            I => \N__21851\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__21879\,
            I => \N__21851\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__21874\,
            I => \N__21851\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21851\
        );

    \I__5278\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21848\
        );

    \I__5277\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21845\
        );

    \I__5276\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21842\
        );

    \I__5275\ : Span4Mux_s2_v
    port map (
            O => \N__21863\,
            I => \N__21837\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__21860\,
            I => \N__21837\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__21851\,
            I => \N__21834\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__21848\,
            I => \N__21831\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21828\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21825\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__21837\,
            I => \N__21822\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__21834\,
            I => \N__21819\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__21831\,
            I => \N__21816\
        );

    \I__5266\ : Span4Mux_s2_v
    port map (
            O => \N__21828\,
            I => \N__21813\
        );

    \I__5265\ : Span4Mux_s2_v
    port map (
            O => \N__21825\,
            I => \N__21810\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__21822\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__21819\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__21816\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__21813\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__21810\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__5259\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__5257\ : Span4Mux_s1_h
    port map (
            O => \N__21793\,
            I => \N__21788\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__21792\,
            I => \N__21785\
        );

    \I__5255\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21777\
        );

    \I__5254\ : Span4Mux_h
    port map (
            O => \N__21788\,
            I => \N__21770\
        );

    \I__5253\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21761\
        );

    \I__5252\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21761\
        );

    \I__5251\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21761\
        );

    \I__5250\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21761\
        );

    \I__5249\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21756\
        );

    \I__5248\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21756\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__21777\,
            I => \N__21753\
        );

    \I__5246\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21744\
        );

    \I__5245\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21744\
        );

    \I__5244\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21744\
        );

    \I__5243\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21744\
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__21770\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__21761\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__21756\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__21753\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__21744\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__21733\,
            I => \N__21730\
        );

    \I__5236\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__21724\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__5233\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__21718\,
            I => \buart.Z_tx.un1_bitcount_c2\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__21715\,
            I => \N__21703\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__21714\,
            I => \N__21699\
        );

    \I__5229\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21679\
        );

    \I__5228\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21679\
        );

    \I__5227\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21679\
        );

    \I__5226\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21679\
        );

    \I__5225\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21679\
        );

    \I__5224\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21679\
        );

    \I__5223\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21679\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21679\
        );

    \I__5221\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21669\
        );

    \I__5220\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21669\
        );

    \I__5219\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21669\
        );

    \I__5218\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21669\
        );

    \I__5217\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21664\
        );

    \I__5216\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21664\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21661\
        );

    \I__5214\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21658\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__21669\,
            I => \N__21654\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__21664\,
            I => \N__21651\
        );

    \I__5211\ : Span4Mux_h
    port map (
            O => \N__21661\,
            I => \N__21648\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__21658\,
            I => \N__21645\
        );

    \I__5209\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21642\
        );

    \I__5208\ : Span12Mux_s3_v
    port map (
            O => \N__21654\,
            I => \N__21639\
        );

    \I__5207\ : Span4Mux_s3_v
    port map (
            O => \N__21651\,
            I => \N__21636\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__21648\,
            I => \N__21631\
        );

    \I__5205\ : Span4Mux_s3_h
    port map (
            O => \N__21645\,
            I => \N__21631\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__21642\,
            I => vbuf_tx_data_rdy
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__21639\,
            I => vbuf_tx_data_rdy
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__21636\,
            I => vbuf_tx_data_rdy
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__21631\,
            I => vbuf_tx_data_rdy
        );

    \I__5200\ : CEMux
    port map (
            O => \N__21622\,
            I => \N__21618\
        );

    \I__5199\ : CEMux
    port map (
            O => \N__21621\,
            I => \N__21615\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21618\,
            I => \N__21612\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21609\
        );

    \I__5196\ : Span4Mux_h
    port map (
            O => \N__21612\,
            I => \N__21606\
        );

    \I__5195\ : Span12Mux_s4_h
    port map (
            O => \N__21609\,
            I => \N__21603\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__21606\,
            I => \N__21600\
        );

    \I__5193\ : Odrv12
    port map (
            O => \N__21603\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__21600\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__5191\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21591\
        );

    \I__5190\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21588\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__21591\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__21588\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__21583\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21566\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21566\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21566\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21566\
        );

    \I__5182\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21561\
        );

    \I__5181\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21561\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21566\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21561\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__5178\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21550\
        );

    \I__5177\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21543\
        );

    \I__5176\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21543\
        );

    \I__5175\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21543\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__21550\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__21543\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21530\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21525\
        );

    \I__5169\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21525\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21530\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__21525\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__21520\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__5165\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21508\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21508\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21501\
        );

    \I__5162\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21501\
        );

    \I__5161\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21501\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__21508\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21501\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__21493\,
            I => \buart.Z_tx.un1_bitcount_c3\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__21490\,
            I => \Lab_UT.dictrl.g0_6_3_cascade_\
        );

    \I__5155\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21481\
        );

    \I__5154\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21481\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21478\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__21475\,
            I => \Lab_UT.dictrl.N_57_0\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21469\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__21469\,
            I => \Lab_UT.dictrl.g0_6_3\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21460\
        );

    \I__5147\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21460\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__21460\,
            I => \Lab_UT.dictrl.g1_1\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__21457\,
            I => \N__21453\
        );

    \I__5144\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21448\
        );

    \I__5143\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21448\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21445\
        );

    \I__5141\ : Odrv12
    port map (
            O => \N__21445\,
            I => \Lab_UT.dictrl.gZ0Z2\
        );

    \I__5140\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21432\
        );

    \I__5139\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21432\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__21440\,
            I => \N__21420\
        );

    \I__5137\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21413\
        );

    \I__5136\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21408\
        );

    \I__5135\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21408\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21405\
        );

    \I__5133\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21402\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21393\
        );

    \I__5131\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21393\
        );

    \I__5130\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21393\
        );

    \I__5129\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21393\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21390\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21387\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21382\
        );

    \I__5125\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21382\
        );

    \I__5124\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21377\
        );

    \I__5123\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21377\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21368\
        );

    \I__5121\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21368\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21365\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__21413\,
            I => \N__21360\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21360\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__21405\,
            I => \N__21344\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21344\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21393\,
            I => \N__21344\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21344\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__21387\,
            I => \N__21344\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21344\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21377\,
            I => \N__21344\
        );

    \I__5110\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21339\
        );

    \I__5109\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21339\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21334\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21334\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21368\,
            I => \N__21329\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21365\,
            I => \N__21329\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__21360\,
            I => \N__21326\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21323\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__21344\,
            I => \N__21318\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__21339\,
            I => \N__21318\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21334\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__21329\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__21326\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21323\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__21318\,
            I => \Lab_UT_dictrl_state_1\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21304\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21300\
        );

    \I__5093\ : InMux
    port map (
            O => \N__21303\,
            I => \N__21297\
        );

    \I__5092\ : Span4Mux_v
    port map (
            O => \N__21300\,
            I => \N__21294\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21297\,
            I => \Lab_UT.dictrl.N_55_0\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__21294\,
            I => \Lab_UT.dictrl.N_55_0\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__21289\,
            I => \N__21284\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21279\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21274\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21271\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21268\
        );

    \I__5084\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21265\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__21279\,
            I => \N__21262\
        );

    \I__5082\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21259\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__21277\,
            I => \N__21256\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21274\,
            I => \N__21252\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21247\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21244\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21265\,
            I => \N__21241\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__21262\,
            I => \N__21236\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__21259\,
            I => \N__21236\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21231\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21231\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__21252\,
            I => \N__21222\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21219\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21216\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__21247\,
            I => \N__21211\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__21244\,
            I => \N__21211\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__21241\,
            I => \N__21204\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__21236\,
            I => \N__21204\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21204\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21195\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21195\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21195\
        );

    \I__5061\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21195\
        );

    \I__5060\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21192\
        );

    \I__5059\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21189\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__21222\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__21219\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__21216\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__21211\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__21204\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21195\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__21192\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__21189\,
            I => \Lab_UT.state_i_4_3\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__21172\,
            I => \Lab_UT.dictrl.g1_rn_0_cascade_\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21160\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21160\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21154\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21154\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21150\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21147\
        );

    \I__5043\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21144\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21136\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21132\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21129\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__21147\,
            I => \N__21126\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21123\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21120\
        );

    \I__5036\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21111\
        );

    \I__5035\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21111\
        );

    \I__5034\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21111\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21111\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__21136\,
            I => \N__21103\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21100\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21097\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__21129\,
            I => \N__21092\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__21126\,
            I => \N__21092\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__21123\,
            I => \N__21085\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21085\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21111\,
            I => \N__21085\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21080\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21080\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21073\
        );

    \I__5021\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21073\
        );

    \I__5020\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21073\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__21103\,
            I => \Lab_UT.state_2\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__21100\,
            I => \Lab_UT.state_2\
        );

    \I__5017\ : Odrv12
    port map (
            O => \N__21097\,
            I => \Lab_UT.state_2\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__21092\,
            I => \Lab_UT.state_2\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__21085\,
            I => \Lab_UT.state_2\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21080\,
            I => \Lab_UT.state_2\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__21073\,
            I => \Lab_UT.state_2\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21055\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21052\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__21052\,
            I => \N__21049\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__21049\,
            I => \N__21046\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__21046\,
            I => \Lab_UT.dictrl.G_25_i_a5_1_0_0\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__21043\,
            I => \N__21037\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__21042\,
            I => \N__21029\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__21041\,
            I => \N__21026\
        );

    \I__5004\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21017\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21014\
        );

    \I__5002\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21011\
        );

    \I__5001\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21008\
        );

    \I__5000\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21005\
        );

    \I__4999\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21002\
        );

    \I__4998\ : InMux
    port map (
            O => \N__21032\,
            I => \N__20999\
        );

    \I__4997\ : InMux
    port map (
            O => \N__21029\,
            I => \N__20994\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21026\,
            I => \N__20994\
        );

    \I__4995\ : InMux
    port map (
            O => \N__21025\,
            I => \N__20989\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21024\,
            I => \N__20989\
        );

    \I__4993\ : InMux
    port map (
            O => \N__21023\,
            I => \N__20986\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21022\,
            I => \N__20983\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21021\,
            I => \N__20978\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21020\,
            I => \N__20978\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__20975\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__20928\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__20925\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__20922\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20919\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20916\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20913\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20910\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__20989\,
            I => \N__20907\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__20986\,
            I => \N__20892\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__20983\,
            I => \N__20889\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20886\
        );

    \I__4977\ : Glb2LocalMux
    port map (
            O => \N__20975\,
            I => \N__20749\
        );

    \I__4976\ : SRMux
    port map (
            O => \N__20974\,
            I => \N__20749\
        );

    \I__4975\ : SRMux
    port map (
            O => \N__20973\,
            I => \N__20749\
        );

    \I__4974\ : SRMux
    port map (
            O => \N__20972\,
            I => \N__20749\
        );

    \I__4973\ : SRMux
    port map (
            O => \N__20971\,
            I => \N__20749\
        );

    \I__4972\ : SRMux
    port map (
            O => \N__20970\,
            I => \N__20749\
        );

    \I__4971\ : SRMux
    port map (
            O => \N__20969\,
            I => \N__20749\
        );

    \I__4970\ : SRMux
    port map (
            O => \N__20968\,
            I => \N__20749\
        );

    \I__4969\ : SRMux
    port map (
            O => \N__20967\,
            I => \N__20749\
        );

    \I__4968\ : SRMux
    port map (
            O => \N__20966\,
            I => \N__20749\
        );

    \I__4967\ : SRMux
    port map (
            O => \N__20965\,
            I => \N__20749\
        );

    \I__4966\ : SRMux
    port map (
            O => \N__20964\,
            I => \N__20749\
        );

    \I__4965\ : SRMux
    port map (
            O => \N__20963\,
            I => \N__20749\
        );

    \I__4964\ : SRMux
    port map (
            O => \N__20962\,
            I => \N__20749\
        );

    \I__4963\ : SRMux
    port map (
            O => \N__20961\,
            I => \N__20749\
        );

    \I__4962\ : SRMux
    port map (
            O => \N__20960\,
            I => \N__20749\
        );

    \I__4961\ : SRMux
    port map (
            O => \N__20959\,
            I => \N__20749\
        );

    \I__4960\ : SRMux
    port map (
            O => \N__20958\,
            I => \N__20749\
        );

    \I__4959\ : SRMux
    port map (
            O => \N__20957\,
            I => \N__20749\
        );

    \I__4958\ : SRMux
    port map (
            O => \N__20956\,
            I => \N__20749\
        );

    \I__4957\ : SRMux
    port map (
            O => \N__20955\,
            I => \N__20749\
        );

    \I__4956\ : SRMux
    port map (
            O => \N__20954\,
            I => \N__20749\
        );

    \I__4955\ : SRMux
    port map (
            O => \N__20953\,
            I => \N__20749\
        );

    \I__4954\ : SRMux
    port map (
            O => \N__20952\,
            I => \N__20749\
        );

    \I__4953\ : SRMux
    port map (
            O => \N__20951\,
            I => \N__20749\
        );

    \I__4952\ : SRMux
    port map (
            O => \N__20950\,
            I => \N__20749\
        );

    \I__4951\ : SRMux
    port map (
            O => \N__20949\,
            I => \N__20749\
        );

    \I__4950\ : SRMux
    port map (
            O => \N__20948\,
            I => \N__20749\
        );

    \I__4949\ : SRMux
    port map (
            O => \N__20947\,
            I => \N__20749\
        );

    \I__4948\ : SRMux
    port map (
            O => \N__20946\,
            I => \N__20749\
        );

    \I__4947\ : SRMux
    port map (
            O => \N__20945\,
            I => \N__20749\
        );

    \I__4946\ : SRMux
    port map (
            O => \N__20944\,
            I => \N__20749\
        );

    \I__4945\ : SRMux
    port map (
            O => \N__20943\,
            I => \N__20749\
        );

    \I__4944\ : SRMux
    port map (
            O => \N__20942\,
            I => \N__20749\
        );

    \I__4943\ : SRMux
    port map (
            O => \N__20941\,
            I => \N__20749\
        );

    \I__4942\ : SRMux
    port map (
            O => \N__20940\,
            I => \N__20749\
        );

    \I__4941\ : SRMux
    port map (
            O => \N__20939\,
            I => \N__20749\
        );

    \I__4940\ : SRMux
    port map (
            O => \N__20938\,
            I => \N__20749\
        );

    \I__4939\ : SRMux
    port map (
            O => \N__20937\,
            I => \N__20749\
        );

    \I__4938\ : SRMux
    port map (
            O => \N__20936\,
            I => \N__20749\
        );

    \I__4937\ : SRMux
    port map (
            O => \N__20935\,
            I => \N__20749\
        );

    \I__4936\ : SRMux
    port map (
            O => \N__20934\,
            I => \N__20749\
        );

    \I__4935\ : SRMux
    port map (
            O => \N__20933\,
            I => \N__20749\
        );

    \I__4934\ : SRMux
    port map (
            O => \N__20932\,
            I => \N__20749\
        );

    \I__4933\ : SRMux
    port map (
            O => \N__20931\,
            I => \N__20749\
        );

    \I__4932\ : Glb2LocalMux
    port map (
            O => \N__20928\,
            I => \N__20749\
        );

    \I__4931\ : Glb2LocalMux
    port map (
            O => \N__20925\,
            I => \N__20749\
        );

    \I__4930\ : Glb2LocalMux
    port map (
            O => \N__20922\,
            I => \N__20749\
        );

    \I__4929\ : Glb2LocalMux
    port map (
            O => \N__20919\,
            I => \N__20749\
        );

    \I__4928\ : Glb2LocalMux
    port map (
            O => \N__20916\,
            I => \N__20749\
        );

    \I__4927\ : Glb2LocalMux
    port map (
            O => \N__20913\,
            I => \N__20749\
        );

    \I__4926\ : Glb2LocalMux
    port map (
            O => \N__20910\,
            I => \N__20749\
        );

    \I__4925\ : Glb2LocalMux
    port map (
            O => \N__20907\,
            I => \N__20749\
        );

    \I__4924\ : SRMux
    port map (
            O => \N__20906\,
            I => \N__20749\
        );

    \I__4923\ : SRMux
    port map (
            O => \N__20905\,
            I => \N__20749\
        );

    \I__4922\ : SRMux
    port map (
            O => \N__20904\,
            I => \N__20749\
        );

    \I__4921\ : SRMux
    port map (
            O => \N__20903\,
            I => \N__20749\
        );

    \I__4920\ : SRMux
    port map (
            O => \N__20902\,
            I => \N__20749\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__20901\,
            I => \N__20749\
        );

    \I__4918\ : SRMux
    port map (
            O => \N__20900\,
            I => \N__20749\
        );

    \I__4917\ : SRMux
    port map (
            O => \N__20899\,
            I => \N__20749\
        );

    \I__4916\ : SRMux
    port map (
            O => \N__20898\,
            I => \N__20749\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__20897\,
            I => \N__20749\
        );

    \I__4914\ : SRMux
    port map (
            O => \N__20896\,
            I => \N__20749\
        );

    \I__4913\ : SRMux
    port map (
            O => \N__20895\,
            I => \N__20749\
        );

    \I__4912\ : Glb2LocalMux
    port map (
            O => \N__20892\,
            I => \N__20749\
        );

    \I__4911\ : Glb2LocalMux
    port map (
            O => \N__20889\,
            I => \N__20749\
        );

    \I__4910\ : Glb2LocalMux
    port map (
            O => \N__20886\,
            I => \N__20749\
        );

    \I__4909\ : GlobalMux
    port map (
            O => \N__20749\,
            I => \N__20746\
        );

    \I__4908\ : gio2CtrlBuf
    port map (
            O => \N__20746\,
            I => rst_g
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__20743\,
            I => \N__20735\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20732\
        );

    \I__4905\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20727\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20727\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20724\
        );

    \I__4902\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20719\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20719\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20716\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20711\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__20724\,
            I => \N__20711\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__20719\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__20716\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__20711\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__4894\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20700\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__20703\,
            I => \N__20697\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__20700\,
            I => \N__20694\
        );

    \I__4891\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20691\
        );

    \I__4890\ : Span4Mux_s1_h
    port map (
            O => \N__20694\,
            I => \N__20688\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__20691\,
            I => \N__20674\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__20688\,
            I => \N__20674\
        );

    \I__4887\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20663\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20663\
        );

    \I__4885\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20663\
        );

    \I__4884\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20663\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20663\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20660\
        );

    \I__4881\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20653\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20653\
        );

    \I__4879\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20653\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__20674\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__20663\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20660\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__20653\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__4871\ : Odrv12
    port map (
            O => \N__20635\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__4870\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20628\
        );

    \I__4869\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20625\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__20628\,
            I => \N__20610\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20625\,
            I => \N__20607\
        );

    \I__4866\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20604\
        );

    \I__4865\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20599\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20599\
        );

    \I__4863\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20596\
        );

    \I__4862\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20587\
        );

    \I__4861\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20587\
        );

    \I__4860\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20587\
        );

    \I__4859\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20587\
        );

    \I__4858\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20584\
        );

    \I__4857\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20579\
        );

    \I__4856\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20574\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20574\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__20610\,
            I => \N__20569\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__20607\,
            I => \N__20569\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20566\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20561\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__20596\,
            I => \N__20561\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20556\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20556\
        );

    \I__4847\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20553\
        );

    \I__4846\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20550\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20579\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20574\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__20569\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__20566\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4841\ : Odrv12
    port map (
            O => \N__20561\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__20556\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__20553\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__20550\,
            I => \Lab_UT.stateZ0Z_0\
        );

    \I__4837\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20527\
        );

    \I__4836\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20527\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__20527\,
            I => \Lab_UT.dictrl.N_59\
        );

    \I__4834\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20512\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20508\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20505\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20518\,
            I => \N__20502\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \N__20499\
        );

    \I__4828\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20495\
        );

    \I__4827\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20491\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20512\,
            I => \N__20488\
        );

    \I__4825\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20484\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20478\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20478\
        );

    \I__4822\ : Span4Mux_v
    port map (
            O => \N__20502\,
            I => \N__20475\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20470\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20470\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20465\
        );

    \I__4818\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20462\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__20491\,
            I => \N__20456\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__20488\,
            I => \N__20453\
        );

    \I__4815\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20449\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20446\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__20483\,
            I => \N__20443\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__20478\,
            I => \N__20438\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__20475\,
            I => \N__20433\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20433\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20430\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20427\
        );

    \I__4807\ : Span12Mux_s11_v
    port map (
            O => \N__20465\,
            I => \N__20422\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20422\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20419\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20460\,
            I => \N__20414\
        );

    \I__4803\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20414\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__20456\,
            I => \N__20411\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__20453\,
            I => \N__20408\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20405\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20400\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__20446\,
            I => \N__20400\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20397\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20392\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20392\
        );

    \I__4794\ : Span4Mux_v
    port map (
            O => \N__20438\,
            I => \N__20383\
        );

    \I__4793\ : Span4Mux_s3_h
    port map (
            O => \N__20433\,
            I => \N__20383\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20430\,
            I => \N__20383\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__20427\,
            I => \N__20383\
        );

    \I__4790\ : Span12Mux_s4_v
    port map (
            O => \N__20422\,
            I => \N__20380\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20419\,
            I => bu_rx_data_3
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__20414\,
            I => bu_rx_data_3
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__20411\,
            I => bu_rx_data_3
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__20408\,
            I => bu_rx_data_3
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20405\,
            I => bu_rx_data_3
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__20400\,
            I => bu_rx_data_3
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__20397\,
            I => bu_rx_data_3
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20392\,
            I => bu_rx_data_3
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__20383\,
            I => bu_rx_data_3
        );

    \I__4780\ : Odrv12
    port map (
            O => \N__20380\,
            I => bu_rx_data_3
        );

    \I__4779\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20353\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20353\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20353\,
            I => \N__20349\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20346\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__20349\,
            I => \Lab_UT.dictrl.N_15_0\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__20346\,
            I => \Lab_UT.dictrl.N_15_0\
        );

    \I__4773\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20331\
        );

    \I__4772\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20331\
        );

    \I__4771\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20327\
        );

    \I__4770\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20322\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20319\
        );

    \I__4768\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20316\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20331\,
            I => \N__20313\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20307\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20304\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20298\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20295\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__20322\,
            I => \N__20292\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20287\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20316\,
            I => \N__20287\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__20313\,
            I => \N__20284\
        );

    \I__4758\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20279\
        );

    \I__4757\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20279\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20276\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__20307\,
            I => \N__20269\
        );

    \I__4754\ : Sp12to4
    port map (
            O => \N__20304\,
            I => \N__20269\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20266\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20263\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__20301\,
            I => \N__20258\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20255\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20248\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__20292\,
            I => \N__20248\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__20287\,
            I => \N__20248\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__20284\,
            I => \N__20241\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20241\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__20276\,
            I => \N__20241\
        );

    \I__4743\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20236\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20236\
        );

    \I__4741\ : Span12Mux_v
    port map (
            O => \N__20269\,
            I => \N__20233\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__20266\,
            I => \N__20230\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20227\
        );

    \I__4738\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20220\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20220\
        );

    \I__4736\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20220\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__20255\,
            I => \N__20213\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__20248\,
            I => \N__20213\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__20241\,
            I => \N__20213\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__20236\,
            I => bu_rx_data_2
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__20233\,
            I => bu_rx_data_2
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__20230\,
            I => bu_rx_data_2
        );

    \I__4729\ : Odrv12
    port map (
            O => \N__20227\,
            I => bu_rx_data_2
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__20220\,
            I => bu_rx_data_2
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__20213\,
            I => bu_rx_data_2
        );

    \I__4726\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20195\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20192\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__20198\,
            I => \N__20188\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20178\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__20192\,
            I => \N__20178\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20174\
        );

    \I__4720\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20171\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20166\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20163\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__20185\,
            I => \N__20159\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20156\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20151\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__20178\,
            I => \N__20148\
        );

    \I__4713\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20145\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__20174\,
            I => \N__20140\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20171\,
            I => \N__20140\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20137\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20134\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20166\,
            I => \N__20131\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20163\,
            I => \N__20128\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__20162\,
            I => \N__20123\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20120\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20117\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20114\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20111\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20151\,
            I => \N__20107\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__20148\,
            I => \N__20100\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20145\,
            I => \N__20100\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__20140\,
            I => \N__20100\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20091\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20091\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__20131\,
            I => \N__20091\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__20128\,
            I => \N__20091\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20086\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20086\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20083\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__20120\,
            I => \N__20080\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__20117\,
            I => \N__20077\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20114\,
            I => \N__20074\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20111\,
            I => \N__20071\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20068\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20107\,
            I => \N__20065\
        );

    \I__4684\ : Span4Mux_h
    port map (
            O => \N__20100\,
            I => \N__20062\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__20091\,
            I => \N__20053\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20086\,
            I => \N__20053\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__20083\,
            I => \N__20053\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__20080\,
            I => \N__20053\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__20077\,
            I => bu_rx_data_1
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__20074\,
            I => bu_rx_data_1
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__20071\,
            I => bu_rx_data_1
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20068\,
            I => bu_rx_data_1
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__20065\,
            I => bu_rx_data_1
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__20062\,
            I => bu_rx_data_1
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__20053\,
            I => bu_rx_data_1
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__20038\,
            I => \N__20034\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20025\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20022\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20019\
        );

    \I__4668\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20016\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20011\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20008\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__20029\,
            I => \N__20004\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__20028\,
            I => \N__20001\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__19998\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__19995\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__20019\,
            I => \N__19992\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20016\,
            I => \N__19987\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20015\,
            I => \N__19982\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19982\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__19977\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__19977\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20007\,
            I => \N__19974\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19969\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19969\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__19998\,
            I => \N__19966\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__19995\,
            I => \N__19961\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__19992\,
            I => \N__19961\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19958\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19955\
        );

    \I__4647\ : Span4Mux_s3_v
    port map (
            O => \N__19987\,
            I => \N__19946\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19946\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__19977\,
            I => \N__19946\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19946\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19969\,
            I => \N__19943\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__19966\,
            I => bu_rx_data_3_rep2
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__19961\,
            I => bu_rx_data_3_rep2
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__19958\,
            I => bu_rx_data_3_rep2
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__19955\,
            I => bu_rx_data_3_rep2
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__19946\,
            I => bu_rx_data_3_rep2
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__19943\,
            I => bu_rx_data_3_rep2
        );

    \I__4636\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__19924\,
            I => \G_6_0_a6_2\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__19921\,
            I => \N__19915\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__19920\,
            I => \N__19912\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__19919\,
            I => \N__19909\
        );

    \I__4630\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19902\
        );

    \I__4629\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19899\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19896\
        );

    \I__4627\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19891\
        );

    \I__4626\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19886\
        );

    \I__4625\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19886\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19881\
        );

    \I__4623\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19881\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__19902\,
            I => \N__19876\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19876\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19873\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19870\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19865\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19852\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19886\,
            I => \N__19852\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19881\,
            I => \N__19852\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__19876\,
            I => \N__19852\
        );

    \I__4613\ : Span4Mux_h
    port map (
            O => \N__19873\,
            I => \N__19852\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19852\
        );

    \I__4611\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19849\
        );

    \I__4610\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19846\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__19865\,
            I => \N__19843\
        );

    \I__4608\ : Span4Mux_v
    port map (
            O => \N__19852\,
            I => \N__19840\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__19849\,
            I => \N__19835\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19846\,
            I => \N__19835\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__19843\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__19840\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4603\ : Odrv12
    port map (
            O => \N__19835\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19811\
        );

    \I__4601\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19811\
        );

    \I__4600\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19808\
        );

    \I__4599\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19801\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19801\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19801\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19795\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19795\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19790\
        );

    \I__4593\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19790\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19783\
        );

    \I__4591\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19783\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19783\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19780\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19773\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__19801\,
            I => \N__19773\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19770\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__19795\,
            I => \N__19767\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19762\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19783\,
            I => \N__19762\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__19780\,
            I => \N__19759\
        );

    \I__4581\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19754\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19754\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__19773\,
            I => \N__19751\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N_63_mux\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__19767\,
            I => \N_63_mux\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__19762\,
            I => \N_63_mux\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__19759\,
            I => \N_63_mux\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__19754\,
            I => \N_63_mux\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__19751\,
            I => \N_63_mux\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19727\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19724\
        );

    \I__4569\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19720\
        );

    \I__4568\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19715\
        );

    \I__4567\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19715\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19710\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19707\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19704\
        );

    \I__4563\ : CascadeMux
    port map (
            O => \N__19723\,
            I => \N__19701\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19696\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19696\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19692\
        );

    \I__4559\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19688\
        );

    \I__4558\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19685\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__19707\,
            I => \N__19680\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__19704\,
            I => \N__19680\
        );

    \I__4555\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19677\
        );

    \I__4554\ : Span4Mux_v
    port map (
            O => \N__19696\,
            I => \N__19674\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19671\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__19692\,
            I => \N__19668\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19665\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__19688\,
            I => \N__19656\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__19685\,
            I => \N__19656\
        );

    \I__4548\ : Span4Mux_v
    port map (
            O => \N__19680\,
            I => \N__19656\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19656\
        );

    \I__4546\ : Span4Mux_s2_v
    port map (
            O => \N__19674\,
            I => \N__19653\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19671\,
            I => \N__19646\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__19668\,
            I => \N__19646\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19646\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__19656\,
            I => \N__19643\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__19653\,
            I => bu_rx_data_3_rep1
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__19646\,
            I => bu_rx_data_3_rep1
        );

    \I__4539\ : Odrv4
    port map (
            O => \N__19643\,
            I => bu_rx_data_3_rep1
        );

    \I__4538\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19633\,
            I => \N__19628\
        );

    \I__4536\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19624\
        );

    \I__4535\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19621\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__19628\,
            I => \N__19618\
        );

    \I__4533\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19615\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__19624\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__19621\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__19618\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__19615\,
            I => \Lab_UT.dictrl.N_72_mux\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19603\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19603\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__19600\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19591\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19591\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19584\
        );

    \I__4522\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19579\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19579\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19575\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19572\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__19584\,
            I => \N__19567\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19567\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19564\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19575\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19572\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__19567\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19564\,
            I => \Lab_UT.dictrl.m13_out\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19552\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19552\,
            I => \N__19549\
        );

    \I__4509\ : Odrv12
    port map (
            O => \N__19549\,
            I => \Lab_UT.dictrl.N_59_1_0\
        );

    \I__4508\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19541\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__19545\,
            I => \N__19538\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__19544\,
            I => \N__19535\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19532\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19529\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19526\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__19532\,
            I => \N__19523\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19518\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__19526\,
            I => \N__19518\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__19523\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__4498\ : Odrv12
    port map (
            O => \N__19518\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__4497\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19509\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19506\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19509\,
            I => \N__19503\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__19506\,
            I => bu_rx_data_fast_0
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__19503\,
            I => bu_rx_data_fast_0
        );

    \I__4492\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19495\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__19495\,
            I => \N__19491\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__19494\,
            I => \N__19488\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__19491\,
            I => \N__19485\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19482\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__19485\,
            I => bu_rx_data_fast_7
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__19482\,
            I => bu_rx_data_fast_7
        );

    \I__4485\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__4483\ : Span4Mux_s3_h
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__19468\,
            I => \Lab_UT.dictrl.g1_1Z0Z_5\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19461\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19458\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19446\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19446\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19443\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19438\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19438\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19435\
        );

    \I__4473\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19430\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19430\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19427\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__19446\,
            I => \N__19420\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19443\,
            I => \N__19420\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19420\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19435\,
            I => \N__19417\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19430\,
            I => bu_rx_data_1_rep1
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19427\,
            I => bu_rx_data_1_rep1
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__19420\,
            I => bu_rx_data_1_rep1
        );

    \I__4463\ : Odrv12
    port map (
            O => \N__19417\,
            I => bu_rx_data_1_rep1
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \Lab_UT.dictrl.g1_1_4_cascade_\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__19405\,
            I => \N__19400\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19395\
        );

    \I__4459\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19392\
        );

    \I__4458\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19385\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19385\
        );

    \I__4456\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19385\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__19395\,
            I => bu_rx_data_6_rep1
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19392\,
            I => bu_rx_data_6_rep1
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__19385\,
            I => bu_rx_data_6_rep1
        );

    \I__4452\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19375\,
            I => \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19357\
        );

    \I__4446\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19352\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19352\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__19360\,
            I => bu_rx_data_5_rep1
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__19357\,
            I => bu_rx_data_5_rep1
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19352\,
            I => bu_rx_data_5_rep1
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__19345\,
            I => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_\
        );

    \I__4440\ : CEMux
    port map (
            O => \N__19342\,
            I => \N__19338\
        );

    \I__4439\ : CEMux
    port map (
            O => \N__19341\,
            I => \N__19335\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19332\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19335\,
            I => \N__19328\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__19332\,
            I => \N__19324\
        );

    \I__4435\ : CEMux
    port map (
            O => \N__19331\,
            I => \N__19321\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__19328\,
            I => \N__19318\
        );

    \I__4433\ : CEMux
    port map (
            O => \N__19327\,
            I => \N__19315\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__19324\,
            I => \N__19310\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19310\
        );

    \I__4430\ : Span4Mux_s2_h
    port map (
            O => \N__19318\,
            I => \N__19307\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19315\,
            I => \N__19304\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__19310\,
            I => \N__19301\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__19307\,
            I => \Lab_UT.g0_0\
        );

    \I__4426\ : Odrv12
    port map (
            O => \N__19304\,
            I => \Lab_UT.g0_0\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__19301\,
            I => \Lab_UT.g0_0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19287\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19284\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__19287\,
            I => \N__19281\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19284\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__19281\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__19276\,
            I => \N__19271\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__19275\,
            I => \N__19268\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__19274\,
            I => \N__19260\
        );

    \I__4415\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19247\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19247\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19247\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19247\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19239\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19239\
        );

    \I__4409\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19232\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19232\
        );

    \I__4407\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19232\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19219\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19219\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19219\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19216\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19213\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__19245\,
            I => \N__19210\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19205\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19239\,
            I => \N__19202\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19199\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19231\,
            I => \N__19192\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19192\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19192\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19187\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19187\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19184\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__19219\,
            I => \N__19181\
        );

    \I__4390\ : Span4Mux_v
    port map (
            O => \N__19216\,
            I => \N__19176\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19213\,
            I => \N__19176\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19173\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19168\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19168\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19161\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__19202\,
            I => \N__19161\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__19199\,
            I => \N__19161\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19158\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19187\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19184\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__19181\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__19176\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__19173\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19168\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__19161\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4374\ : Odrv12
    port map (
            O => \N__19158\,
            I => \Lab_UT.un1_next_state66_0\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__19141\,
            I => \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19132\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19132\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__19129\,
            I => \N__19126\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__19126\,
            I => \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19118\
        );

    \I__4366\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19113\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19113\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19107\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19107\
        );

    \I__4362\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19104\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__19107\,
            I => \N__19101\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19104\,
            I => m7_a0
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__19101\,
            I => m7_a0
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__19096\,
            I => \Lab_UT.dictrl.N_8_0_cascade_\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__19093\,
            I => \Lab_UT.dictrl.G_6_0_0_1_cascade_\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19087\,
            I => \Lab_UT.dictrl.G_6_0_0\
        );

    \I__4354\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__19081\,
            I => \Lab_UT.dictrl.N_8_0\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19075\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__19075\,
            I => \Lab_UT.dictrl.i9_mux\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__19072\,
            I => \N__19065\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__19071\,
            I => \N__19058\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19055\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19042\
        );

    \I__4346\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19042\
        );

    \I__4345\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19042\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19035\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19035\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19035\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19031\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19027\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19055\,
            I => \N__19024\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19021\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19018\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19015\
        );

    \I__4335\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19008\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19008\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19008\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19003\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19003\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19000\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19031\,
            I => \N__18997\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19030\,
            I => \N__18994\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__18989\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__19024\,
            I => \N__18989\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19021\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19018\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__19015\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19008\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__19003\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19000\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__18997\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18994\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4317\ : Odrv4
    port map (
            O => \N__18989\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__18970\,
            I => \N__18966\
        );

    \I__4315\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18962\
        );

    \I__4314\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18957\
        );

    \I__4313\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18957\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__18962\,
            I => \Lab_UT.dictrl.N_60\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__18957\,
            I => \Lab_UT.dictrl.N_60\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__18952\,
            I => \Lab_UT.dictrl.i8_mux_cascade_\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__18949\,
            I => \N__18945\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18942\
        );

    \I__4307\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18939\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__18942\,
            I => \N__18932\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__18939\,
            I => \N__18929\
        );

    \I__4304\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18924\
        );

    \I__4303\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18924\
        );

    \I__4302\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18921\
        );

    \I__4301\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18917\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__18932\,
            I => \N__18914\
        );

    \I__4299\ : Span4Mux_h
    port map (
            O => \N__18929\,
            I => \N__18907\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18907\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18907\
        );

    \I__4296\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18904\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__18917\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__18914\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__18907\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__18904\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__4291\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18892\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__18892\,
            I => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__18889\,
            I => \Lab_UT.dictrl.m34_0_cascade_\
        );

    \I__4288\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18883\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__18883\,
            I => \N__18880\
        );

    \I__4286\ : Span4Mux_v
    port map (
            O => \N__18880\,
            I => \N__18875\
        );

    \I__4285\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18870\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18870\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__18875\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18870\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__18865\,
            I => \Lab_UT.dictrl.next_state_1_3_cascade_\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__18862\,
            I => \N__18858\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__18861\,
            I => \N__18854\
        );

    \I__4278\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18847\
        );

    \I__4277\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18847\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18847\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__18844\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__4273\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__4272\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18835\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18832\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__18832\,
            I => \Lab_UT.dictrl.N_33_0\
        );

    \I__4269\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__18826\,
            I => \N__18823\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__18823\,
            I => \Lab_UT.dictrl.N_60_0_0\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__18820\,
            I => \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18805\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18805\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18805\
        );

    \I__4262\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18805\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18805\,
            I => \Lab_UT.dictrl.N_26_0\
        );

    \I__4260\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18796\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18796\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__18793\,
            I => \N__18790\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__18790\,
            I => \Lab_UT.dictrl.i8_mux_0\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18781\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18781\,
            I => \Lab_UT.dictrl.m34_0\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18774\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18771\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__18774\,
            I => \N__18764\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__18771\,
            I => \N__18764\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__18770\,
            I => \N__18761\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__18769\,
            I => \N__18758\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__18764\,
            I => \N__18755\
        );

    \I__4245\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18750\
        );

    \I__4244\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18750\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__18755\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18750\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__18745\,
            I => \N__18742\
        );

    \I__4240\ : InMux
    port map (
            O => \N__18742\,
            I => \N__18737\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__18741\,
            I => \N__18734\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \N__18730\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18727\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18723\
        );

    \I__4235\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18718\
        );

    \I__4234\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18718\
        );

    \I__4233\ : Span4Mux_h
    port map (
            O => \N__18727\,
            I => \N__18715\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18726\,
            I => \N__18712\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__18723\,
            I => \N__18709\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__18718\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__18715\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18712\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4227\ : Odrv12
    port map (
            O => \N__18709\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__18700\,
            I => \N__18696\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18690\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18690\
        );

    \I__4223\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18687\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18690\,
            I => \N__18684\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18681\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__18684\,
            I => \N__18678\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__18681\,
            I => \N__18675\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__18678\,
            I => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__18675\,
            I => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18667\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__18667\,
            I => \Lab_UT.dictrl.g0_1_mb_rn_0\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__18664\,
            I => \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18661\,
            I => \N__18658\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__18658\,
            I => \N__18654\
        );

    \I__4211\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18651\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__18654\,
            I => \N__18648\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18645\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__18648\,
            I => \N__18642\
        );

    \I__4207\ : Span4Mux_h
    port map (
            O => \N__18645\,
            I => \N__18639\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__18642\,
            I => \Lab_UT.dictrl.N_57_1\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__18639\,
            I => \Lab_UT.dictrl.N_57_1\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18627\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__18630\,
            I => \N__18624\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18621\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18618\
        );

    \I__4199\ : Span4Mux_s3_v
    port map (
            O => \N__18621\,
            I => \N__18615\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18618\,
            I => \N__18612\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__18615\,
            I => \N__18607\
        );

    \I__4196\ : Span4Mux_s3_h
    port map (
            O => \N__18612\,
            I => \N__18607\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__18607\,
            I => \N__18604\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__18604\,
            I => \Lab_UT.dictrl.N_55_1\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18594\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18597\,
            I => \N__18590\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18594\,
            I => \N__18587\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18582\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18582\
        );

    \I__4187\ : Span4Mux_v
    port map (
            O => \N__18587\,
            I => \N__18579\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__18582\,
            I => \N__18576\
        );

    \I__4185\ : Span4Mux_v
    port map (
            O => \N__18579\,
            I => \N__18573\
        );

    \I__4184\ : Span4Mux_v
    port map (
            O => \N__18576\,
            I => \N__18570\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__18573\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__18570\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__18565\,
            I => \Lab_UT.dictrl.next_state_1_2_cascade_\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18552\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18552\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18552\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__18559\,
            I => \N__18549\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18552\,
            I => \N__18546\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__18546\,
            I => \Lab_UT.dictrl.state_i_4_2\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18543\,
            I => \Lab_UT.dictrl.state_i_4_2\
        );

    \I__4172\ : CEMux
    port map (
            O => \N__18538\,
            I => \N__18534\
        );

    \I__4171\ : CEMux
    port map (
            O => \N__18537\,
            I => \N__18531\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18534\,
            I => \N__18527\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18531\,
            I => \N__18523\
        );

    \I__4168\ : CEMux
    port map (
            O => \N__18530\,
            I => \N__18520\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__18527\,
            I => \N__18517\
        );

    \I__4166\ : CEMux
    port map (
            O => \N__18526\,
            I => \N__18514\
        );

    \I__4165\ : Span4Mux_s3_h
    port map (
            O => \N__18523\,
            I => \N__18509\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__18520\,
            I => \N__18509\
        );

    \I__4163\ : Sp12to4
    port map (
            O => \N__18517\,
            I => \N__18506\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18514\,
            I => \N__18501\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__18509\,
            I => \N__18501\
        );

    \I__4160\ : Odrv12
    port map (
            O => \N__18506\,
            I => \Lab_UT.bu_rx_data_rdy_0\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__18501\,
            I => \Lab_UT.bu_rx_data_rdy_0\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18490\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18495\,
            I => \N__18490\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18490\,
            I => \Lab_UT.dictrl.g0_1_mb_sn\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18483\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18479\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__18483\,
            I => \N__18476\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18473\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18479\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__18476\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18473\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__18466\,
            I => \Lab_UT.dictrl.un15_loadalarm_0_cascade_\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18460\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__18460\,
            I => \Lab_UT.dictrl.loadalarm_0_0\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18452\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__18456\,
            I => \N__18449\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__18455\,
            I => \N__18444\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18452\,
            I => \N__18441\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18438\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__18448\,
            I => \N__18435\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18447\,
            I => \N__18429\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18423\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__18441\,
            I => \N__18418\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__18438\,
            I => \N__18418\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18412\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18405\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18405\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18405\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18429\,
            I => \N__18402\
        );

    \I__4130\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18395\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18395\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18395\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18423\,
            I => \N__18390\
        );

    \I__4126\ : Span4Mux_h
    port map (
            O => \N__18418\,
            I => \N__18390\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18417\,
            I => \N__18383\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18383\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18383\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18412\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18405\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__18402\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18395\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__18390\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__18383\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18365\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18351\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18351\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18346\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18341\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18341\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18332\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18332\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18332\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18332\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18327\
        );

    \I__4105\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18327\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18321\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18351\,
            I => \N__18316\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18311\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18311\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__18346\,
            I => \N__18308\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__18341\,
            I => \N__18301\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18332\,
            I => \N__18301\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18301\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18294\
        );

    \I__4095\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18294\
        );

    \I__4094\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18294\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18321\,
            I => \N__18291\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18286\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18286\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__18316\,
            I => \N__18283\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18311\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__18308\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__18301\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__18294\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__18291\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__18286\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__18283\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18253\
        );

    \I__4080\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18253\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18253\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18249\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__18261\,
            I => \N__18245\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18239\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18253\,
            I => \N__18236\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18233\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18230\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18227\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18222\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18222\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18217\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18217\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18239\,
            I => \N__18213\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__18236\,
            I => \N__18208\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__18233\,
            I => \N__18208\
        );

    \I__4064\ : Span4Mux_v
    port map (
            O => \N__18230\,
            I => \N__18203\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18203\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18198\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18198\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18195\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__18213\,
            I => \N__18192\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__18208\,
            I => \N__18189\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__18203\,
            I => \N__18186\
        );

    \I__4056\ : Span12Mux_s8_h
    port map (
            O => \N__18198\,
            I => \N__18183\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__18195\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__18192\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__18189\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__18186\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__4051\ : Odrv12
    port map (
            O => \N__18183\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18160\
        );

    \I__4049\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18160\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18160\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18160\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__18160\,
            I => \N__18154\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18150\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18158\,
            I => \N__18147\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18144\
        );

    \I__4042\ : Span4Mux_s3_h
    port map (
            O => \N__18154\,
            I => \N__18141\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18138\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18150\,
            I => \N__18133\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18133\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18144\,
            I => \Lab_UT.next_state_1\
        );

    \I__4037\ : Odrv4
    port map (
            O => \N__18141\,
            I => \Lab_UT.next_state_1\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18138\,
            I => \Lab_UT.next_state_1\
        );

    \I__4035\ : Odrv12
    port map (
            O => \N__18133\,
            I => \Lab_UT.next_state_1\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18115\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18106\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18106\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18106\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18106\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18119\,
            I => \N__18103\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18100\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18097\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18106\,
            I => \Lab_UT.next_state_2\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__18103\,
            I => \Lab_UT.next_state_2\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18100\,
            I => \Lab_UT.next_state_2\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__18097\,
            I => \Lab_UT.next_state_2\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__18088\,
            I => \N__18084\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__18087\,
            I => \N__18080\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18075\
        );

    \I__4019\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18068\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18068\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18068\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18062\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__18075\,
            I => \N__18057\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18057\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18050\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18050\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18050\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18047\
        );

    \I__4009\ : Span4Mux_v
    port map (
            O => \N__18057\,
            I => \N__18041\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18041\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__18047\,
            I => \N__18037\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18034\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__18041\,
            I => \N__18031\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18028\
        );

    \I__4003\ : Sp12to4
    port map (
            O => \N__18037\,
            I => \N__18023\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__18034\,
            I => \N__18023\
        );

    \I__4001\ : Span4Mux_h
    port map (
            O => \N__18031\,
            I => \N__18020\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18028\,
            I => bu_rx_data_rdy
        );

    \I__3999\ : Odrv12
    port map (
            O => \N__18023\,
            I => bu_rx_data_rdy
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__18020\,
            I => bu_rx_data_rdy
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__18013\,
            I => \N__18008\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18012\,
            I => \N__18005\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__18011\,
            I => \N__18002\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18008\,
            I => \N__17999\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__17996\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17993\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__17999\,
            I => \N__17989\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__17996\,
            I => \N__17984\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17984\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17981\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__17989\,
            I => \N__17978\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__17984\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__17981\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__17978\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \Lab_UT.didp.countrce3.q_5_1_cascade_\
        );

    \I__3982\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17961\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17958\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__17961\,
            I => \N__17953\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__17958\,
            I => \N__17953\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__17953\,
            I => \N__17949\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17946\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__17949\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__17946\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17937\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__17940\,
            I => \N__17934\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17926\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17923\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17920\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17913\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17913\
        );

    \I__3966\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17913\
        );

    \I__3965\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17910\
        );

    \I__3964\ : Span4Mux_v
    port map (
            O => \N__17926\,
            I => \N__17905\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17923\,
            I => \N__17905\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17920\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17913\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__17910\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__17905\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__17896\,
            I => \N__17891\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \N__17886\
        );

    \I__3956\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17881\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17881\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17878\
        );

    \I__3953\ : InMux
    port map (
            O => \N__17889\,
            I => \N__17873\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17873\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__17881\,
            I => \N__17870\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17866\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17863\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__17870\,
            I => \N__17860\
        );

    \I__3947\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17857\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__17866\,
            I => \N__17854\
        );

    \I__3945\ : Span12Mux_s8_h
    port map (
            O => \N__17863\,
            I => \N__17851\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__17860\,
            I => \N__17848\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__17857\,
            I => \N__17843\
        );

    \I__3942\ : Span4Mux_s2_v
    port map (
            O => \N__17854\,
            I => \N__17843\
        );

    \I__3941\ : Odrv12
    port map (
            O => \N__17851\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__17848\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__17843\,
            I => \Lab_UT.state_ret_8_ess\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__17836\,
            I => \N__17832\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__17835\,
            I => \N__17828\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17815\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17815\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17815\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17815\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17810\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17810\
        );

    \I__3930\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17806\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17803\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__17810\,
            I => \N__17800\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17797\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17806\,
            I => \Lab_UT.next_state_0\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__17803\,
            I => \Lab_UT.next_state_0\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__17800\,
            I => \Lab_UT.next_state_0\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17797\,
            I => \Lab_UT.next_state_0\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17785\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17782\
        );

    \I__3920\ : Odrv12
    port map (
            O => \N__17782\,
            I => \Lab_UT.didp.N_90\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17779\,
            I => \N__17776\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__17776\,
            I => \N__17773\
        );

    \I__3917\ : Odrv12
    port map (
            O => \N__17773\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17767\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17767\,
            I => \Lab_UT.LdSones_i_4\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__17764\,
            I => \N__17759\
        );

    \I__3913\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17756\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17753\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17750\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__17756\,
            I => \N__17747\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17739\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17750\,
            I => \N__17739\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__17747\,
            I => \N__17739\
        );

    \I__3906\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17736\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__17739\,
            I => \N__17733\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17736\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__17733\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__3902\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17722\
        );

    \I__3901\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17718\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17714\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17711\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__17722\,
            I => \N__17708\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17705\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__17718\,
            I => \N__17702\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17699\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17696\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17693\
        );

    \I__3892\ : Span4Mux_h
    port map (
            O => \N__17708\,
            I => \N__17690\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17681\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__17702\,
            I => \N__17681\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17699\,
            I => \N__17681\
        );

    \I__3888\ : Span4Mux_h
    port map (
            O => \N__17696\,
            I => \N__17678\
        );

    \I__3887\ : Span4Mux_s2_v
    port map (
            O => \N__17693\,
            I => \N__17675\
        );

    \I__3886\ : Span4Mux_v
    port map (
            O => \N__17690\,
            I => \N__17672\
        );

    \I__3885\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17667\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17667\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__17681\,
            I => \N__17664\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__17678\,
            I => \N__17659\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__17675\,
            I => \N__17659\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__17672\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__17667\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__17664\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__17659\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17647\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17643\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17640\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__17643\,
            I => \N__17635\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__17640\,
            I => \N__17632\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17629\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \N__17626\
        );

    \I__3869\ : Span4Mux_h
    port map (
            O => \N__17635\,
            I => \N__17623\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__17632\,
            I => \N__17620\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17629\,
            I => \N__17617\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17626\,
            I => \N__17614\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__17623\,
            I => \Lab_UT.LdSones\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__17620\,
            I => \Lab_UT.LdSones\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__17617\,
            I => \Lab_UT.LdSones\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__17614\,
            I => \Lab_UT.LdSones\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17595\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17595\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17595\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17592\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__17595\,
            I => \N__17586\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__17592\,
            I => \N__17583\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17579\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17575\
        );

    \I__3853\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17572\
        );

    \I__3852\ : Span4Mux_h
    port map (
            O => \N__17586\,
            I => \N__17569\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__17583\,
            I => \N__17566\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17563\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17579\,
            I => \N__17560\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17557\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17575\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17572\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__17569\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__17566\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17563\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__17560\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17557\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3840\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__17536\,
            I => \Lab_UT.didp.countrce1.q_5_1\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__17533\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17527\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17527\,
            I => \Lab_UT.didp.countrce3.q_5_3\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17524\,
            I => \Lab_UT.didp.countrce1.un13_qPone_cascade_\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17511\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17511\
        );

    \I__3831\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17511\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17496\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17493\
        );

    \I__3828\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17490\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17479\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17479\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17479\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17479\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17479\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17470\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17470\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17470\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17470\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17467\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17464\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17461\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__17493\,
            I => \N__17456\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17456\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17451\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17470\,
            I => \N__17451\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17467\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17464\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__17461\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__17456\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__17451\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17434\
        );

    \I__3804\ : Span4Mux_h
    port map (
            O => \N__17434\,
            I => \N__17426\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17423\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17418\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17418\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17415\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17412\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__17426\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17423\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17418\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17415\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17412\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17393\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17390\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17387\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__17393\,
            I => \N__17384\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17390\,
            I => \N__17381\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17387\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__17384\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3785\ : Odrv12
    port map (
            O => \N__17381\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17368\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__17373\,
            I => \N__17364\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__17372\,
            I => \N__17360\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__17371\,
            I => \N__17356\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17368\,
            I => \N__17353\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17340\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17340\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17340\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17340\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17340\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17356\,
            I => \N__17340\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__17353\,
            I => \N__17337\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17334\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__17337\,
            I => \Lab_UT.min1_2\
        );

    \I__3770\ : Odrv12
    port map (
            O => \N__17334\,
            I => \Lab_UT.min1_2\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17326\,
            I => \Lab_UT.didp.countrce1.q_5_2\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__17323\,
            I => \N__17320\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17316\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__17319\,
            I => \N__17313\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17309\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17306\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17303\
        );

    \I__3761\ : Sp12to4
    port map (
            O => \N__17309\,
            I => \N__17297\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17306\,
            I => \N__17297\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17294\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17291\
        );

    \I__3757\ : Span12Mux_s6_h
    port map (
            O => \N__17297\,
            I => \N__17286\
        );

    \I__3756\ : Span12Mux_s5_h
    port map (
            O => \N__17294\,
            I => \N__17286\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17283\
        );

    \I__3754\ : Odrv12
    port map (
            O => \N__17286\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__17283\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17272\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17277\,
            I => \N__17272\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17263\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17259\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17256\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__17266\,
            I => \N__17253\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__17263\,
            I => \N__17250\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17247\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17259\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17256\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__17253\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__17250\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17247\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17232\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17228\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17232\,
            I => \N__17222\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17219\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__17228\,
            I => \N__17216\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17213\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17208\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17208\
        );

    \I__3730\ : Span4Mux_h
    port map (
            O => \N__17222\,
            I => \N__17205\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17202\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__17216\,
            I => \N__17197\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17197\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17208\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__17205\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3724\ : Odrv12
    port map (
            O => \N__17202\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__17197\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17184\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__17187\,
            I => \N__17181\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17184\,
            I => \N__17177\
        );

    \I__3719\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17172\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__17180\,
            I => \N__17169\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__17177\,
            I => \N__17166\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17163\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17160\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17157\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17154\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__17166\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17163\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17160\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17157\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17154\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17134\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17134\
        );

    \I__3705\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17134\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__17134\,
            I => \N__17131\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__17131\,
            I => \N__17128\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__17128\,
            I => \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__3700\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17118\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17114\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__17118\,
            I => \N__17111\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17105\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17114\,
            I => \N__17102\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__17111\,
            I => \N__17099\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17094\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17094\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17091\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17105\,
            I => \N__17088\
        );

    \I__3690\ : Sp12to4
    port map (
            O => \N__17102\,
            I => \N__17081\
        );

    \I__3689\ : Sp12to4
    port map (
            O => \N__17099\,
            I => \N__17081\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17081\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17078\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__17088\,
            I => \N__17075\
        );

    \I__3685\ : Span12Mux_s5_h
    port map (
            O => \N__17081\,
            I => \N__17072\
        );

    \I__3684\ : Span12Mux_v
    port map (
            O => \N__17078\,
            I => \N__17069\
        );

    \I__3683\ : Span4Mux_v
    port map (
            O => \N__17075\,
            I => \N__17066\
        );

    \I__3682\ : Odrv12
    port map (
            O => \N__17072\,
            I => \Lab_UT.LdMtens\
        );

    \I__3681\ : Odrv12
    port map (
            O => \N__17069\,
            I => \Lab_UT.LdMtens\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__17066\,
            I => \Lab_UT.LdMtens\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17053\,
            I => \Lab_UT.didp.countrce4.un20_qPone\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__17047\,
            I => \N__17041\
        );

    \I__3674\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17037\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17034\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17031\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__17041\,
            I => \N__17028\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17025\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17037\,
            I => \N__17022\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17034\,
            I => \N__17019\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__17031\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__17028\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17025\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__17022\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__17019\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17008\,
            I => \N__17005\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17005\,
            I => \Lab_UT.didp.countrce4.q_5_3\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16997\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16989\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16989\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16986\
        );

    \I__3656\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16982\
        );

    \I__3655\ : InMux
    port map (
            O => \N__16995\,
            I => \N__16977\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16977\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16974\
        );

    \I__3652\ : Span4Mux_h
    port map (
            O => \N__16986\,
            I => \N__16971\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16968\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__16982\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__16977\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3648\ : Odrv12
    port map (
            O => \N__16974\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__16971\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16968\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16950\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16945\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16945\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16942\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__16953\,
            I => \N__16938\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__16950\,
            I => \N__16931\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16931\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__16942\,
            I => \N__16931\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16928\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16925\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__16931\,
            I => \N__16922\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16919\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__16925\,
            I => \Lab_UT.LdMones\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__16922\,
            I => \Lab_UT.LdMones\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__16919\,
            I => \Lab_UT.LdMones\
        );

    \I__3630\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16901\
        );

    \I__3629\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16901\
        );

    \I__3628\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16890\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16890\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16890\
        );

    \I__3625\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16890\
        );

    \I__3624\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16890\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__16901\,
            I => \Lab_UT.sec2_0\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16890\,
            I => \Lab_UT.sec2_0\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__16885\,
            I => \N__16878\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__16884\,
            I => \N__16875\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__16883\,
            I => \N__16871\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__16882\,
            I => \N__16867\
        );

    \I__3617\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16862\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16862\
        );

    \I__3615\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16851\
        );

    \I__3614\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16851\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16851\
        );

    \I__3612\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16851\
        );

    \I__3611\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16851\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__16862\,
            I => \Lab_UT.sec2_3\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__16851\,
            I => \Lab_UT.sec2_3\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__16846\,
            I => \N__16841\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__16845\,
            I => \N__16837\
        );

    \I__3606\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16823\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16823\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16823\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16823\
        );

    \I__3602\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16823\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16818\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16818\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16815\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__16818\,
            I => \Lab_UT.sec2_1\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__16815\,
            I => \Lab_UT.sec2_1\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__16810\,
            I => \N__16807\
        );

    \I__3595\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16796\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16796\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16785\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16785\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16803\,
            I => \N__16785\
        );

    \I__3590\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16785\
        );

    \I__3589\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16785\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__16796\,
            I => \Lab_UT.sec2_2\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__16785\,
            I => \Lab_UT.sec2_2\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16776\
        );

    \I__3585\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16773\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16776\,
            I => \N__16770\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__16773\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3582\ : Odrv12
    port map (
            O => \N__16770\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3581\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16756\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16753\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16750\
        );

    \I__3577\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16747\
        );

    \I__3576\ : Span4Mux_h
    port map (
            O => \N__16756\,
            I => \N__16744\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__16753\,
            I => \N__16739\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16739\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16747\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__16744\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__16739\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16726\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__16720\,
            I => \uu2.bitmap_RNIM5E21Z0Z_314\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16710\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16703\
        );

    \I__3563\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16703\
        );

    \I__3562\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16703\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16700\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__16710\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__16703\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16700\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16690\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16684\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__16684\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16678\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__16678\,
            I => \uu2.N_152\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16672\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16672\,
            I => \N__16668\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16665\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__16668\,
            I => \N__16662\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__16665\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__16662\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16651\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16651\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16651\,
            I => \N__16647\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16644\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__16647\,
            I => \N__16639\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__16644\,
            I => \N__16639\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__16639\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16628\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16625\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \N__16621\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16614\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16614\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16614\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16628\,
            I => \N__16611\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16608\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16605\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16602\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16614\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__16611\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__16608\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16605\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16602\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16587\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16583\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__16587\,
            I => \N__16580\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16586\,
            I => \N__16577\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__16583\,
            I => \N__16574\
        );

    \I__3518\ : Span4Mux_v
    port map (
            O => \N__16580\,
            I => \N__16569\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__16577\,
            I => \N__16569\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__16574\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__16569\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16561\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__16561\,
            I => \N__16552\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16539\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16539\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16539\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16539\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16539\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16539\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__16552\,
            I => \N__16536\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16539\,
            I => \N__16533\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__16536\,
            I => \Lab_UT.min1_1\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__16533\,
            I => \Lab_UT.min1_1\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__16528\,
            I => \N__16525\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16522\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__16522\,
            I => \Lab_UT.didp.countrce4.un13_qPone\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16516\,
            I => \Lab_UT.didp.countrce4.q_5_2\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16510\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16510\,
            I => \N__16507\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__16507\,
            I => \N__16504\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__16504\,
            I => \uu2.bitmap_pmux_20_ns_1\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16498\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__16495\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16489\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16489\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16483\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__16483\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16477\
        );

    \I__3485\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16474\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16471\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__16471\,
            I => \uu2.bitmap_pmux_26_bm_1\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__16468\,
            I => \N__16464\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__16467\,
            I => \N__16459\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16464\,
            I => \N__16454\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16451\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16446\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16446\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16441\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16441\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__16454\,
            I => \N__16436\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16436\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__16446\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__16441\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3470\ : Odrv12
    port map (
            O => \N__16436\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16426\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__16423\,
            I => \uu2.bitmap_RNIP2JO1Z0Z_34\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16411\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16398\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16398\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16398\
        );

    \I__3462\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16398\
        );

    \I__3461\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16398\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16398\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16395\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__16398\,
            I => \Lab_UT.min1_0\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__16395\,
            I => \Lab_UT.min1_0\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__16390\,
            I => \N__16384\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__16389\,
            I => \N__16380\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16376\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__16387\,
            I => \N__16372\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16359\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16359\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16359\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16359\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16359\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16359\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16356\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16353\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16356\,
            I => \N__16350\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__16353\,
            I => \Lab_UT.min1_3\
        );

    \I__3442\ : Odrv12
    port map (
            O => \N__16350\,
            I => \Lab_UT.min1_3\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16342\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__16342\,
            I => \N__16339\
        );

    \I__3439\ : Span4Mux_h
    port map (
            O => \N__16339\,
            I => \N__16336\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__16336\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16326\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16332\,
            I => \N__16326\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16318\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16326\,
            I => \N__16315\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \N__16312\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16306\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16323\,
            I => \N__16299\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16299\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16299\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__16318\,
            I => \N__16294\
        );

    \I__3427\ : Span4Mux_v
    port map (
            O => \N__16315\,
            I => \N__16294\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16289\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16289\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16286\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16283\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__16306\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16299\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__16294\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16289\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__16286\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16283\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16267\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16264\,
            I => \N__16259\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16263\,
            I => \N__16256\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__16262\,
            I => \N__16252\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16246\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16237\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16237\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16237\
        );

    \I__3407\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16237\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16250\,
            I => \N__16231\
        );

    \I__3405\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16228\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__16246\,
            I => \N__16223\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16223\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16216\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16216\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16216\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16213\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16228\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__16223\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__16216\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__16213\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16201\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16195\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__16195\,
            I => \N__16192\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__16192\,
            I => \uu2.bitmap_pmux_19_ns_1\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16182\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16177\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16177\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16172\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16172\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16167\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16167\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16172\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__16167\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__16162\,
            I => \uu2.un3_w_addr_user_4_cascade_\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16156\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16156\,
            I => \uu2.un3_w_addr_user_5\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16147\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16147\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16147\,
            I => \N__16144\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__16144\,
            I => \N__16141\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__16141\,
            I => \uu2.un3_w_addr_user\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16137\,
            I => \N__16129\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__16136\,
            I => \N__16123\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__16135\,
            I => \N__16120\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16116\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16129\,
            I => \N__16113\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16128\,
            I => \N__16108\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16103\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16103\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16098\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16098\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16095\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__16116\,
            I => \N__16092\
        );

    \I__3359\ : Span4Mux_s1_v
    port map (
            O => \N__16113\,
            I => \N__16089\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16112\,
            I => \N__16084\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16084\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16081\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__16103\,
            I => \N__16072\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16072\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16095\,
            I => \N__16072\
        );

    \I__3352\ : Span4Mux_s1_v
    port map (
            O => \N__16092\,
            I => \N__16072\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__16089\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16084\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16081\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__16072\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__16063\,
            I => \N__16060\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__3344\ : Odrv12
    port map (
            O => \N__16054\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16044\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16041\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16036\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16036\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16033\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16044\,
            I => \N__16026\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16026\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16026\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16033\,
            I => \N__16023\
        );

    \I__3334\ : Odrv12
    port map (
            O => \N__16026\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__16023\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \N__16015\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__3330\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16004\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16004\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16001\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__16009\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16004\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__16001\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__15994\,
            I => \N__15990\
        );

    \I__3323\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15979\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15979\
        );

    \I__3321\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15979\
        );

    \I__3320\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15979\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15979\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15973\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__15970\,
            I => \N__15963\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15954\
        );

    \I__3314\ : InMux
    port map (
            O => \N__15968\,
            I => \N__15954\
        );

    \I__3313\ : InMux
    port map (
            O => \N__15967\,
            I => \N__15954\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15966\,
            I => \N__15951\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__15963\,
            I => \N__15948\
        );

    \I__3310\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15943\
        );

    \I__3309\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15943\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__15954\,
            I => \N__15940\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__15951\,
            I => \N__15935\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__15948\,
            I => \N__15935\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15943\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__15940\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__15935\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \N__15924\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15916\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15916\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15916\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15916\,
            I => \N__15912\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15909\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__15912\,
            I => \uu2.un404_ci\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__15909\,
            I => \uu2.un404_ci\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \N__15899\
        );

    \I__3293\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15894\
        );

    \I__3292\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15894\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15891\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__15894\,
            I => \N__15888\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__15891\,
            I => \N__15885\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__15888\,
            I => \uu2.un426_ci_3\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__15885\,
            I => \uu2.un426_ci_3\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \uu2.un404_ci_cascade_\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15874\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__15874\,
            I => \uu2.vbuf_w_addr_user.un448_ci_0\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15868\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15863\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15858\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15858\
        );

    \I__3279\ : Odrv12
    port map (
            O => \N__15863\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__15858\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__3277\ : CEMux
    port map (
            O => \N__15853\,
            I => \N__15850\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__15850\,
            I => \N__15847\
        );

    \I__3275\ : Sp12to4
    port map (
            O => \N__15847\,
            I => \N__15844\
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__15844\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__3273\ : SRMux
    port map (
            O => \N__15841\,
            I => \N__15838\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15835\
        );

    \I__3271\ : Span4Mux_s0_v
    port map (
            O => \N__15835\,
            I => \N__15831\
        );

    \I__3270\ : SRMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__15831\,
            I => \N__15823\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15823\
        );

    \I__3267\ : Span4Mux_s0_v
    port map (
            O => \N__15823\,
            I => \N__15819\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15816\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15819\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_4\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15816\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_4\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15808\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15808\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15802\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15802\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__15799\,
            I => \N__15796\
        );

    \I__3258\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15790\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15790\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15790\,
            I => \N__15780\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15775\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15775\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__15787\,
            I => \N__15772\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15769\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__15785\,
            I => \N__15766\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__15784\,
            I => \N__15762\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15759\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__15780\,
            I => \N__15754\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15775\,
            I => \N__15754\
        );

    \I__3246\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15751\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__15769\,
            I => \N__15748\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15745\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15740\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15740\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15759\,
            I => \N__15737\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__15754\,
            I => \N__15734\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15727\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__15748\,
            I => \N__15727\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15727\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__15740\,
            I => \N__15724\
        );

    \I__3235\ : Odrv12
    port map (
            O => \N__15737\,
            I => bu_rx_data_2_rep1
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__15734\,
            I => bu_rx_data_2_rep1
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__15727\,
            I => bu_rx_data_2_rep1
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__15724\,
            I => bu_rx_data_2_rep1
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15705\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15700\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15700\
        );

    \I__3227\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15695\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15692\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15705\,
            I => \N__15687\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15687\
        );

    \I__3223\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15682\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15682\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__15695\,
            I => \N__15679\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15676\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__15687\,
            I => \N__15673\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15682\,
            I => \N__15670\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__15679\,
            I => bu_rx_data_0_rep1
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__15676\,
            I => bu_rx_data_0_rep1
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__15673\,
            I => bu_rx_data_0_rep1
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__15670\,
            I => bu_rx_data_0_rep1
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15661\,
            I => \N__15658\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15655\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15655\,
            I => \N__15652\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__15652\,
            I => \G_6_0_a6_3_3\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15649\,
            I => \N__15642\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15648\,
            I => \N__15637\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15637\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15632\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15645\,
            I => \N__15632\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__15642\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15637\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15632\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15618\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15615\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15606\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15606\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15606\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15606\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15615\,
            I => bu_rx_data_7_rep1
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15606\,
            I => bu_rx_data_7_rep1
        );

    \I__3193\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15594\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15594\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15591\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15594\,
            I => \N__15586\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__15591\,
            I => \N__15586\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__15586\,
            I => \N__15582\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15585\,
            I => \N__15579\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__3184\ : Span4Mux_v
    port map (
            O => \N__15576\,
            I => \N__15568\
        );

    \I__3183\ : Span4Mux_s3_v
    port map (
            O => \N__15573\,
            I => \N__15568\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__15568\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__15565\,
            I => \N__15555\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15550\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15547\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15544\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15541\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15536\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15536\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15533\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15526\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15526\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15526\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15550\,
            I => \N__15521\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15547\,
            I => \N__15512\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15544\,
            I => \N__15512\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15512\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15536\,
            I => \N__15512\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__15533\,
            I => \N__15507\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15526\,
            I => \N__15507\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15504\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15501\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__15521\,
            I => \N__15498\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__15512\,
            I => \N__15495\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__15507\,
            I => \N__15492\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__15504\,
            I => bu_rx_data_7
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15501\,
            I => bu_rx_data_7
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__15498\,
            I => bu_rx_data_7
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__15495\,
            I => bu_rx_data_7
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__15492\,
            I => bu_rx_data_7
        );

    \I__3153\ : CEMux
    port map (
            O => \N__15481\,
            I => \N__15454\
        );

    \I__3152\ : CEMux
    port map (
            O => \N__15480\,
            I => \N__15454\
        );

    \I__3151\ : CEMux
    port map (
            O => \N__15479\,
            I => \N__15454\
        );

    \I__3150\ : CEMux
    port map (
            O => \N__15478\,
            I => \N__15454\
        );

    \I__3149\ : CEMux
    port map (
            O => \N__15477\,
            I => \N__15454\
        );

    \I__3148\ : CEMux
    port map (
            O => \N__15476\,
            I => \N__15454\
        );

    \I__3147\ : CEMux
    port map (
            O => \N__15475\,
            I => \N__15454\
        );

    \I__3146\ : CEMux
    port map (
            O => \N__15474\,
            I => \N__15454\
        );

    \I__3145\ : CEMux
    port map (
            O => \N__15473\,
            I => \N__15454\
        );

    \I__3144\ : GlobalMux
    port map (
            O => \N__15454\,
            I => \N__15451\
        );

    \I__3143\ : gio2CtrlBuf
    port map (
            O => \N__15451\,
            I => \buart.Z_rx.sample_g\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \N__15445\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15440\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15444\,
            I => \N__15434\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15434\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15431\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15428\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15434\,
            I => \N__15425\
        );

    \I__3135\ : Span4Mux_h
    port map (
            O => \N__15431\,
            I => \N__15422\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15428\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__15425\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__15422\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__15415\,
            I => \Lab_UT.dictrl.m22_xZ0Z1_cascade_\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \Lab_UT.dictrl.N_72_mux_cascade_\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15406\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15397\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15394\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15391\
        );

    \I__3124\ : Span4Mux_s3_v
    port map (
            O => \N__15400\,
            I => \N__15379\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__15397\,
            I => \N__15379\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__15394\,
            I => \N__15372\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__15391\,
            I => \N__15372\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15369\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15366\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15361\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15361\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15354\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15354\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15354\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__15379\,
            I => \N__15351\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15346\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15346\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__15372\,
            I => bu_rx_data_4
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15369\,
            I => bu_rx_data_4
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15366\,
            I => bu_rx_data_4
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15361\,
            I => bu_rx_data_4
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__15354\,
            I => bu_rx_data_4
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__15351\,
            I => bu_rx_data_4
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15346\,
            I => bu_rx_data_4
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__15331\,
            I => \N__15328\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15324\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \N__15321\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15318\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__15318\,
            I => \N__15312\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15315\,
            I => bu_rx_data_fast_3
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__15312\,
            I => bu_rx_data_fast_3
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__15307\,
            I => \N__15303\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__15306\,
            I => \N__15300\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15303\,
            I => \N__15294\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15291\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__15291\,
            I => \N__15285\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__15288\,
            I => \Lab_UT.dictrl.m34Z0Z_1\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__15285\,
            I => \Lab_UT.dictrl.m34Z0Z_1\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \Lab_UT.dictrl.g1_0_xZ0Z1_cascade_\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15274\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15274\,
            I => \N__15271\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__15271\,
            I => \Lab_UT.dictrl.g1_0_4\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15265\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15265\,
            I => \Lab_UT.dictrl.g0_5_3\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__15262\,
            I => \Lab_UT.dictrl.g1_0_cascade_\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15252\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15252\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15249\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15252\,
            I => \N__15245\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15249\,
            I => \N__15242\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15239\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__15245\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15242\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__15239\,
            I => \Lab_UT.dictrl.m22Z0Z_4\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15229\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__15229\,
            I => \Lab_UT.dictrl.g0_5Z0Z_4\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15220\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15215\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15215\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15212\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15220\,
            I => \N__15207\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15207\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__15212\,
            I => \N__15202\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__15207\,
            I => \N__15202\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__15202\,
            I => \Lab_UT.dictrl.next_state66_2\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__15199\,
            I => \N__15195\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15198\,
            I => \N__15191\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15188\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15180\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15177\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15174\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15169\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15169\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15162\
        );

    \I__3050\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15162\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15162\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15180\,
            I => \N__15159\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15152\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__15174\,
            I => \N__15152\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15169\,
            I => \N__15152\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15162\,
            I => \N__15149\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__15159\,
            I => \N__15146\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__15152\,
            I => \N__15143\
        );

    \I__3041\ : Sp12to4
    port map (
            O => \N__15149\,
            I => \N__15140\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__15146\,
            I => \Lab_UT.dictrl.state_i_3_0\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__15143\,
            I => \Lab_UT.dictrl.state_i_3_0\
        );

    \I__3038\ : Odrv12
    port map (
            O => \N__15140\,
            I => \Lab_UT.dictrl.state_i_3_0\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__15133\,
            I => \N_5_cascade_\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15130\,
            I => \N__15127\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15127\,
            I => \N__15124\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__15124\,
            I => \N__15121\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__15121\,
            I => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__15118\,
            I => \Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15111\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15108\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15111\,
            I => \Lab_UT.dictrl.N_67_mux\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15108\,
            I => \Lab_UT.dictrl.N_67_mux\
        );

    \I__3027\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__15100\,
            I => \N__15097\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__15097\,
            I => \Lab_UT.dictrl.G_6_0_1_0\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15091\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15091\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__3022\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15082\
        );

    \I__3021\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15082\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15079\
        );

    \I__3019\ : Odrv12
    port map (
            O => \N__15079\,
            I => \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15073\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15073\,
            I => \Lab_UT.dictrl.g0_3_4\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15067\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__15067\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15061\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__15058\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__15058\,
            I => \Lab_UT.dictrl.G_14_0_a2_4_2\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__15055\,
            I => \N__15051\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15054\,
            I => \N__15048\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15037\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15037\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15037\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15037\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__15034\,
            I => \Lab_UT.dictrl.G_14_0_0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15031\,
            I => \N__15028\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15025\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__15025\,
            I => \Lab_UT.dictrl.g2_0_0\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__15022\,
            I => \N__15019\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15016\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15016\,
            I => \shifter_1_rep1_RNI0FPF\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15010\,
            I => \N__14998\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15009\,
            I => \N__14998\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15008\,
            I => \N__14998\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15007\,
            I => \N__14998\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__14998\,
            I => \N__14995\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__14995\,
            I => \Lab_UT.dictrl.G_14_0_1\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14989\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N_15\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__14986\,
            I => \Lab_UT.dictrl.G_14_0_a2_1_cascade_\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14977\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14977\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14977\,
            I => \N_14_0\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__14974\,
            I => \N__14968\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__14973\,
            I => \N__14965\
        );

    \I__2982\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14956\
        );

    \I__2981\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14956\
        );

    \I__2980\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14956\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14956\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__14956\,
            I => \N__14953\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__14953\,
            I => \N__14950\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__14950\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__14947\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_\
        );

    \I__2974\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14940\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14943\,
            I => \N__14937\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14940\,
            I => \Lab_UT.dictrl.N_22\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__14937\,
            I => \Lab_UT.dictrl.N_22\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__14932\,
            I => \N__14929\
        );

    \I__2969\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14926\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__14926\,
            I => \Lab_UT.dictrl.next_state_0_1\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__14923\,
            I => \Lab_UT.dictrl.N_20_0_0_cascade_\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14917\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__14917\,
            I => \Lab_UT.dictrl.N_22_0_0\
        );

    \I__2964\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14911\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14911\,
            I => \Lab_UT.didp.g0_0Z0Z_2\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__14908\,
            I => \Lab_UT.next_state_1_0_0_1_cascade_\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14899\
        );

    \I__2960\ : InMux
    port map (
            O => \N__14904\,
            I => \N__14899\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__14899\,
            I => \N__14896\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__14896\,
            I => \Lab_UT.dictrl.next_state6\
        );

    \I__2957\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__2956\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14887\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__14887\,
            I => \Lab_UT.dictrl.m19_1\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__14884\,
            I => \N__14881\
        );

    \I__2953\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14878\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14875\
        );

    \I__2951\ : Odrv12
    port map (
            O => \N__14875\,
            I => \Lab_UT.dictrl.m19_1_0\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14868\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__14871\,
            I => \N__14864\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__14868\,
            I => \N__14861\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14858\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14855\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__14861\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14858\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14855\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2942\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__14845\,
            I => \N__14840\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14837\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14834\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__14840\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14837\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__14834\,
            I => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__14827\,
            I => \Lab_UT.dictrl.N_20_cascade_\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14817\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14814\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14817\,
            I => \Lab_UT.dictrl.dicRun_1\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14814\,
            I => \Lab_UT.dictrl.dicRun_1\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14805\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14802\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__14805\,
            I => \Lab_UT.LdASones\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14802\,
            I => \Lab_UT.LdASones\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14794\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14791\
        );

    \I__2923\ : Span4Mux_s3_h
    port map (
            O => \N__14791\,
            I => \N__14787\
        );

    \I__2922\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__14787\,
            I => \N__14781\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14784\,
            I => \N__14778\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__14781\,
            I => \Lab_UT.LdAStens\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__14778\,
            I => \Lab_UT.LdAStens\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14764\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14772\,
            I => \N__14764\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14764\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14761\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__14758\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__14755\,
            I => \N__14751\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__14754\,
            I => \N__14748\
        );

    \I__2909\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14743\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14738\
        );

    \I__2907\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14738\
        );

    \I__2906\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14735\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__14743\,
            I => \N__14732\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14729\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__14735\,
            I => \N__14726\
        );

    \I__2902\ : Span4Mux_h
    port map (
            O => \N__14732\,
            I => \N__14721\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__14729\,
            I => \N__14721\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__14726\,
            I => \N__14718\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__14721\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__14718\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2897\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14707\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14712\,
            I => \N__14707\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__14707\,
            I => \Lab_UT.dictrl.dicLdAMones_1\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14701\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14698\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__14695\,
            I => \Lab_UT.LdAMones\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__14692\,
            I => \Lab_UT.LdAMones_cascade_\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14683\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__14683\,
            I => \N__14680\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__14680\,
            I => \N__14677\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__14677\,
            I => \Lab_UT.dictrl.state_ret_2_fast\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14671\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14659\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14659\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14659\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14654\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14649\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14649\
        );

    \I__2876\ : Span4Mux_s1_v
    port map (
            O => \N__14654\,
            I => \N__14644\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__14649\,
            I => \N__14641\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14636\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14636\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__14644\,
            I => \Lab_UT.min2_2\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__14641\,
            I => \Lab_UT.min2_2\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14636\,
            I => \Lab_UT.min2_2\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__14629\,
            I => \N__14623\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__14628\,
            I => \N__14618\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__14627\,
            I => \N__14615\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14610\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14610\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__14622\,
            I => \N__14606\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14599\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14599\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14599\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__14610\,
            I => \N__14596\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14591\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14591\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14599\,
            I => \Lab_UT.min2_3\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__14596\,
            I => \Lab_UT.min2_3\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__14591\,
            I => \Lab_UT.min2_3\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14578\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14578\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14572\
        );

    \I__2851\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14565\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14565\
        );

    \I__2849\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14565\
        );

    \I__2848\ : Span4Mux_s3_v
    port map (
            O => \N__14572\,
            I => \N__14560\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__14565\,
            I => \N__14557\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14552\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14552\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__14560\,
            I => \Lab_UT.min2_0\
        );

    \I__2843\ : Odrv12
    port map (
            O => \N__14557\,
            I => \Lab_UT.min2_0\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__14552\,
            I => \Lab_UT.min2_0\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__2840\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__14539\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14528\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14525\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14522\
        );

    \I__2834\ : Span4Mux_h
    port map (
            O => \N__14528\,
            I => \N__14517\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14525\,
            I => \N__14517\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14514\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__14517\,
            I => \N__14511\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__14514\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__14511\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14492\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14492\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14492\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__14500\,
            I => \N__14489\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__14499\,
            I => \N__14485\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14492\,
            I => \N__14481\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14476\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14476\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14471\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14471\
        );

    \I__2817\ : Span4Mux_s1_v
    port map (
            O => \N__14481\,
            I => \N__14468\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14476\,
            I => \N__14465\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14471\,
            I => \N__14462\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__14468\,
            I => \Lab_UT.min2_1\
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__14465\,
            I => \Lab_UT.min2_1\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__14462\,
            I => \Lab_UT.min2_1\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__14455\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14445\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14445\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14442\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14445\,
            I => \N__14439\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14434\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__14439\,
            I => \N__14429\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14426\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14423\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__14434\,
            I => \N__14420\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14415\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14415\
        );

    \I__2799\ : Span4Mux_s2_v
    port map (
            O => \N__14429\,
            I => \N__14412\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14426\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14423\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__14420\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14415\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__14412\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14397\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14400\,
            I => \N__14393\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14397\,
            I => \N__14390\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14396\,
            I => \N__14387\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14393\,
            I => \N__14384\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__14390\,
            I => \N__14379\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__14387\,
            I => \N__14379\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__14384\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__14379\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14368\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__14368\,
            I => \N__14365\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__14365\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14359\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14359\,
            I => \N__14354\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14351\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14348\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__14354\,
            I => \N__14344\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14351\,
            I => \N__14339\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14348\,
            I => \N__14339\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14336\
        );

    \I__2772\ : Span4Mux_h
    port map (
            O => \N__14344\,
            I => \N__14333\
        );

    \I__2771\ : Odrv12
    port map (
            O => \N__14339\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__14336\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__14333\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14326\,
            I => \N__14323\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14323\,
            I => \N__14319\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14322\,
            I => \N__14316\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__14319\,
            I => \N__14311\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__14316\,
            I => \N__14311\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__14308\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__14305\,
            I => \N__14302\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14293\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14290\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14285\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14285\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14278\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14278\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14278\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14275\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14290\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14285\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14278\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2749\ : Odrv12
    port map (
            O => \N__14275\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14261\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14254\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14250\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__14261\,
            I => \N__14247\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14244\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14241\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14238\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14235\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14254\,
            I => \N__14232\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14229\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14224\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__14247\,
            I => \N__14224\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14244\,
            I => \N__14216\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14211\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14238\,
            I => \N__14211\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14235\,
            I => \N__14206\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__14232\,
            I => \N__14206\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14229\,
            I => \N__14201\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__14224\,
            I => \N__14201\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14196\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14196\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14189\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14189\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14189\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__14216\,
            I => \N__14186\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__14211\,
            I => \N__14183\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__14206\,
            I => \N__14178\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__14201\,
            I => \N__14178\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__14196\,
            I => \N__14173\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14189\,
            I => \N__14173\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__14186\,
            I => bu_rx_data_0
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__14183\,
            I => bu_rx_data_0
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__14178\,
            I => bu_rx_data_0
        );

    \I__2715\ : Odrv12
    port map (
            O => \N__14173\,
            I => bu_rx_data_0
        );

    \I__2714\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14161\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14161\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14150\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14147\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14144\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__14150\,
            I => \N__14139\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__14147\,
            I => \N__14139\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__14144\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__14139\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__14134\,
            I => \N__14127\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__14133\,
            I => \N__14124\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \N__14121\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14131\,
            I => \N__14118\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14113\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14100\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14100\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14100\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14100\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14100\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14100\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14113\,
            I => \Lab_UT.sec1_1\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14100\,
            I => \Lab_UT.sec1_1\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14086\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14073\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14073\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14073\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14073\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14073\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14073\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__14086\,
            I => \Lab_UT.sec1_2\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14073\,
            I => \Lab_UT.sec1_2\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__14068\,
            I => \N__14059\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__14067\,
            I => \N__14056\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__14066\,
            I => \N__14053\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14065\,
            I => \N__14040\
        );

    \I__2678\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14040\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14040\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14040\
        );

    \I__2675\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14040\
        );

    \I__2674\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14040\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14037\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__14040\,
            I => \N__14034\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14037\,
            I => \Lab_UT.sec1_3\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__14034\,
            I => \Lab_UT.sec1_3\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14020\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14007\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14007\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14007\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14007\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14007\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14007\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__14020\,
            I => \Lab_UT.sec1_0\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__14007\,
            I => \Lab_UT.sec1_0\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13999\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__13999\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13993\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__13993\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13987\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__13987\,
            I => \uu2.bitmap_pmux_17_ns_1\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13979\
        );

    \I__2653\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13972\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13972\
        );

    \I__2651\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13972\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13972\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2649\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13963\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__13963\,
            I => \uu2.bitmap_pmux_16_ns_1\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2645\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13948\
        );

    \I__2644\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13948\
        );

    \I__2643\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13936\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13936\
        );

    \I__2641\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13936\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__13948\,
            I => \N__13933\
        );

    \I__2639\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13925\
        );

    \I__2638\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13925\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13925\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13920\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13920\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__13936\,
            I => \N__13917\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__13933\,
            I => \N__13914\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13911\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__13925\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13920\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__13917\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__13914\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__13911\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13893\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13890\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__13893\,
            I => \N__13885\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__13890\,
            I => \N__13885\
        );

    \I__2621\ : Span4Mux_h
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__13882\,
            I => \uu2.N_44\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__13879\,
            I => \N__13875\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13872\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13868\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13872\,
            I => \N__13865\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13862\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13868\,
            I => \N__13859\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__13865\,
            I => \N__13856\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13862\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__13859\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__13856\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2609\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13846\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__13846\,
            I => \N__13843\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__13843\,
            I => \N__13840\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__13840\,
            I => \Lab_UT.didp.reset_12_1_3\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13834\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__13834\,
            I => \N__13831\
        );

    \I__2603\ : Span4Mux_v
    port map (
            O => \N__13831\,
            I => \N__13828\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__13828\,
            I => \N__13823\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13818\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13818\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__13823\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13818\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13810\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13810\,
            I => \N__13806\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13803\
        );

    \I__2594\ : Span4Mux_s3_v
    port map (
            O => \N__13806\,
            I => \N__13800\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13803\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__13800\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__13789\,
            I => \N__13786\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__13786\,
            I => \N__13781\
        );

    \I__2587\ : InMux
    port map (
            O => \N__13785\,
            I => \N__13778\
        );

    \I__2586\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13775\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__13781\,
            I => \N__13772\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__13778\,
            I => \buart.Z_rx.idle\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__13775\,
            I => \buart.Z_rx.idle\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__13772\,
            I => \buart.Z_rx.idle\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13761\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__13764\,
            I => \N__13754\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13745\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13742\
        );

    \I__2577\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13739\
        );

    \I__2576\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13736\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13733\
        );

    \I__2574\ : InMux
    port map (
            O => \N__13754\,
            I => \N__13730\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13721\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13721\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13721\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13721\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13716\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13716\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__13745\,
            I => \N__13713\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13742\,
            I => \N__13706\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13739\,
            I => \N__13706\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__13736\,
            I => \N__13706\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13703\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__13730\,
            I => \N__13698\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13721\,
            I => \N__13698\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__13716\,
            I => \N__13691\
        );

    \I__2559\ : Span4Mux_s1_h
    port map (
            O => \N__13713\,
            I => \N__13691\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__13706\,
            I => \N__13691\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__13703\,
            I => \N__13686\
        );

    \I__2556\ : Span4Mux_h
    port map (
            O => \N__13698\,
            I => \N__13686\
        );

    \I__2555\ : Sp12to4
    port map (
            O => \N__13691\,
            I => \N__13683\
        );

    \I__2554\ : Sp12to4
    port map (
            O => \N__13686\,
            I => \N__13680\
        );

    \I__2553\ : Span12Mux_s7_h
    port map (
            O => \N__13683\,
            I => \N__13677\
        );

    \I__2552\ : Span12Mux_v
    port map (
            O => \N__13680\,
            I => \N__13674\
        );

    \I__2551\ : Odrv12
    port map (
            O => \N__13677\,
            I => \buart.Z_rx.startbit\
        );

    \I__2550\ : Odrv12
    port map (
            O => \N__13674\,
            I => \buart.Z_rx.startbit\
        );

    \I__2549\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13666\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__13666\,
            I => \N__13663\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__13663\,
            I => \N__13658\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13662\,
            I => \N__13655\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13652\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__13658\,
            I => \N__13649\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13655\,
            I => \N__13646\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13652\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__13649\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__13646\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13639\,
            I => \N__13635\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13632\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13628\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13625\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13622\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__13628\,
            I => \N__13619\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__13625\,
            I => \N__13614\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13614\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__13619\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__13614\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__13609\,
            I => \N__13603\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13596\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13596\
        );

    \I__2526\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13590\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13590\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13585\
        );

    \I__2523\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13585\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13596\,
            I => \N__13582\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13579\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13590\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13585\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__13582\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13579\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13567\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__13567\,
            I => \Lab_UT.didp.countrce2.N_93\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13560\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13555\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13560\,
            I => \N__13552\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13547\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13547\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__13555\,
            I => \N__13543\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__13552\,
            I => \N__13538\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13538\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13535\
        );

    \I__2505\ : Span12Mux_s3_v
    port map (
            O => \N__13543\,
            I => \N__13532\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__13538\,
            I => \N__13529\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13535\,
            I => \o_One_Sec_Pulse\
        );

    \I__2502\ : Odrv12
    port map (
            O => \N__13532\,
            I => \o_One_Sec_Pulse\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__13529\,
            I => \o_One_Sec_Pulse\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13522\,
            I => \N__13519\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13519\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13513\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13513\,
            I => \N__13509\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13512\,
            I => \N__13506\
        );

    \I__2495\ : Span4Mux_s1_v
    port map (
            O => \N__13509\,
            I => \N__13503\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13506\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__13503\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13495\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13495\,
            I => \N__13492\
        );

    \I__2490\ : Span4Mux_s1_v
    port map (
            O => \N__13492\,
            I => \N__13489\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__13489\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13486\,
            I => \N__13483\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13480\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13480\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13474\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13474\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13471\,
            I => \N__13465\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13455\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13455\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13455\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13465\,
            I => \N__13452\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__13464\,
            I => \N__13449\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13446\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13462\,
            I => \N__13443\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13455\,
            I => \N__13438\
        );

    \I__2474\ : Span4Mux_h
    port map (
            O => \N__13452\,
            I => \N__13438\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13435\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13446\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13443\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__13438\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__13435\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__2468\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13421\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13418\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13415\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13421\,
            I => \N__13412\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13418\,
            I => \N__13409\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13415\,
            I => \N__13406\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__13412\,
            I => \N__13403\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__13409\,
            I => \N__13400\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__13406\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__13403\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__13400\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13388\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13392\,
            I => \N__13383\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13383\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__13388\,
            I => \N__13380\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13383\,
            I => \N__13375\
        );

    \I__2452\ : Span12Mux_s6_h
    port map (
            O => \N__13380\,
            I => \N__13375\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__13375\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13372\,
            I => \N__13368\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13365\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13362\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13358\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__13362\,
            I => \N__13355\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13352\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__13358\,
            I => \N__13349\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__13355\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__13352\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__13349\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13333\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13333\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13330\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13327\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13322\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13333\,
            I => \N__13319\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13316\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__13327\,
            I => \N__13313\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__13326\,
            I => \N__13307\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13304\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13322\,
            I => \N__13301\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__13319\,
            I => \N__13298\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__13316\,
            I => \N__13295\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__13313\,
            I => \N__13292\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13283\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13311\,
            I => \N__13283\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13283\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13283\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13304\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__13301\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__13298\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__13295\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__13292\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13283\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__13270\,
            I => \N__13267\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13264\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__13264\,
            I => \uu2.N_45\
        );

    \I__2413\ : CEMux
    port map (
            O => \N__13261\,
            I => \N__13257\
        );

    \I__2412\ : CEMux
    port map (
            O => \N__13260\,
            I => \N__13254\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13250\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__13254\,
            I => \N__13247\
        );

    \I__2409\ : CEMux
    port map (
            O => \N__13253\,
            I => \N__13244\
        );

    \I__2408\ : Span4Mux_s3_v
    port map (
            O => \N__13250\,
            I => \N__13241\
        );

    \I__2407\ : Span4Mux_s0_v
    port map (
            O => \N__13247\,
            I => \N__13238\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13244\,
            I => \N__13233\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__13241\,
            I => \N__13233\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__13238\,
            I => \uu2.N_33_1\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__13233\,
            I => \uu2.N_33_1\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__13225\,
            I => \N__13221\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__13224\,
            I => \N__13216\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__13221\,
            I => \N__13211\
        );

    \I__2398\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13204\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13204\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13204\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13199\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13199\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__13211\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13204\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__13199\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__13192\,
            I => \N__13189\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13189\,
            I => \N__13186\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__13183\,
            I => \N__13180\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__13180\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13167\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13176\,
            I => \N__13164\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13175\,
            I => \N__13161\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13152\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13152\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13152\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13147\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13170\,
            I => \N__13147\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13167\,
            I => \N__13142\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13164\,
            I => \N__13142\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13161\,
            I => \N__13139\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13134\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13134\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__13152\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13147\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__13142\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__13139\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13134\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__13123\,
            I => \N__13120\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13117\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13117\,
            I => \N__13114\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__13114\,
            I => \N__13111\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__13111\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13105\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13105\,
            I => \N__13096\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13091\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13091\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13082\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13082\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13082\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13082\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__13096\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__13091\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__13082\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__13075\,
            I => \N__13072\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13072\,
            I => \N__13069\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13066\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__13066\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__13063\,
            I => \N__13060\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13057\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13057\,
            I => \N__13054\
        );

    \I__2344\ : Odrv12
    port map (
            O => \N__13054\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__13051\,
            I => \Lab_UT.dictrl.g0_3_3_cascade_\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13045\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13045\,
            I => \N__13042\
        );

    \I__2340\ : Odrv12
    port map (
            O => \N__13042\,
            I => \Lab_UT.dictrl.N_72_mux_0\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13035\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13032\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13035\,
            I => \N__13029\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__13032\,
            I => \N__13025\
        );

    \I__2335\ : Span4Mux_h
    port map (
            O => \N__13029\,
            I => \N__13019\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13028\,
            I => \N__13016\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__13025\,
            I => \N__13013\
        );

    \I__2332\ : InMux
    port map (
            O => \N__13024\,
            I => \N__13008\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13008\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13005\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__13019\,
            I => bu_rx_data_fast_2
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13016\,
            I => bu_rx_data_fast_2
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__13013\,
            I => bu_rx_data_fast_2
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13008\,
            I => bu_rx_data_fast_2
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__13005\,
            I => bu_rx_data_fast_2
        );

    \I__2324\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12987\
        );

    \I__2323\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12984\
        );

    \I__2322\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12981\
        );

    \I__2321\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12978\
        );

    \I__2320\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12975\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12987\,
            I => bu_rx_data_fast_1
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__12984\,
            I => bu_rx_data_fast_1
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__12981\,
            I => bu_rx_data_fast_1
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__12978\,
            I => bu_rx_data_fast_1
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12975\,
            I => bu_rx_data_fast_1
        );

    \I__2314\ : InMux
    port map (
            O => \N__12964\,
            I => \N__12959\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12953\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12946\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__12959\,
            I => \N__12943\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12938\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12938\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__12956\,
            I => \N__12934\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__12953\,
            I => \N__12930\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12925\
        );

    \I__2305\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12925\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12920\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12920\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12913\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__12943\,
            I => \N__12913\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__12938\,
            I => \N__12913\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12906\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12906\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12906\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__12930\,
            I => bu_rx_data_6
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__12925\,
            I => bu_rx_data_6
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12920\,
            I => bu_rx_data_6
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__12913\,
            I => bu_rx_data_6
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12906\,
            I => bu_rx_data_6
        );

    \I__2291\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12890\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12894\,
            I => \N__12887\
        );

    \I__2289\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12880\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12890\,
            I => \N__12875\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12887\,
            I => \N__12875\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12872\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12869\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12861\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12858\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__12880\,
            I => \N__12851\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__12875\,
            I => \N__12851\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__12872\,
            I => \N__12851\
        );

    \I__2279\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12844\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12844\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12844\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12837\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12865\,
            I => \N__12837\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12864\,
            I => \N__12837\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12861\,
            I => bu_rx_data_5
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12858\,
            I => bu_rx_data_5
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__12851\,
            I => bu_rx_data_5
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__12844\,
            I => bu_rx_data_5
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12837\,
            I => bu_rx_data_5
        );

    \I__2268\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12822\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12819\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12822\,
            I => \N__12816\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__12819\,
            I => bu_rx_data_fast_6
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__12816\,
            I => bu_rx_data_fast_6
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__12811\,
            I => \N__12805\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12797\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12797\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12797\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12791\
        );

    \I__2258\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12791\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12788\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12785\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12791\,
            I => \N__12780\
        );

    \I__2254\ : Span12Mux_v
    port map (
            O => \N__12788\,
            I => \N__12780\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__12785\,
            I => \uu2.N_40\
        );

    \I__2252\ : Odrv12
    port map (
            O => \N__12780\,
            I => \uu2.N_40\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__12775\,
            I => \Lab_UT.i8_mux_0_cascade_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12769\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12766\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__12766\,
            I => \Lab_UT.didp.g0_0_2Z0Z_1\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12763\,
            I => \N__12760\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12760\,
            I => \Lab_UT.dictrl.g0_0_sn\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__12757\,
            I => \Lab_UT.dictrl.g1_1_0_1_cascade_\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12751\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12751\,
            I => \Lab_UT.g1\
        );

    \I__2242\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12745\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12745\,
            I => \Lab_UT.dictrl.g0_0_rn_0\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__12742\,
            I => \N__12737\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12734\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12729\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12729\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12734\,
            I => \Lab_UT.dictrl.m22Z0Z_1\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12729\,
            I => \Lab_UT.dictrl.m22Z0Z_1\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12719\
        );

    \I__2233\ : IoInMux
    port map (
            O => \N__12723\,
            I => \N__12716\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12712\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12719\,
            I => \N__12709\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__12716\,
            I => \N__12706\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12703\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12712\,
            I => \N__12700\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__12709\,
            I => \N__12697\
        );

    \I__2226\ : IoSpan4Mux
    port map (
            O => \N__12706\,
            I => \N__12694\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12703\,
            I => \N__12691\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__12700\,
            I => \N__12688\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__12697\,
            I => \N__12683\
        );

    \I__2222\ : Span4Mux_s1_h
    port map (
            O => \N__12694\,
            I => \N__12683\
        );

    \I__2221\ : Odrv12
    port map (
            O => \N__12691\,
            I => rst
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__12688\,
            I => rst
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__12683\,
            I => rst
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__12676\,
            I => \Lab_UT.dictrl.g1_1_0_0_cascade_\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12670\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12670\,
            I => \Lab_UT.dictrl.g1_1_0\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12664\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__12664\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12658\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12658\,
            I => \Lab_UT.dictrl.N_3\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__12655\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12649\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12649\,
            I => \Lab_UT.dictrl.m37_N_2LZ0Z1\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12643\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__12643\,
            I => \Lab_UT.dictrl.N_72_mux_1\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__12640\,
            I => \Lab_UT.dictrl.G_25_i_1_cascade_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12634\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12634\,
            I => \Lab_UT.dictrl.G_25_i_0\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12628\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__12628\,
            I => \Lab_UT.dictrl.G_25_i_a5_1_0\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__12625\,
            I => \Lab_UT.dictrl.N_18_0_0_cascade_\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12619\,
            I => \Lab_UT.dictrl.g0_6_3_0\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__12616\,
            I => \N__12613\
        );

    \I__2197\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12610\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__2195\ : Odrv12
    port map (
            O => \N__12607\,
            I => \Lab_UT.dictrl.g2Z0Z_0\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__12604\,
            I => \N__12600\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12596\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12593\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12590\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12596\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12593\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12590\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__12583\,
            I => \Lab_UT.dispString.N_118_cascade_\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12577\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_1\
        );

    \I__2184\ : CEMux
    port map (
            O => \N__12574\,
            I => \N__12571\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__12568\,
            I => \N__12564\
        );

    \I__2181\ : CEMux
    port map (
            O => \N__12567\,
            I => \N__12561\
        );

    \I__2180\ : Span4Mux_v
    port map (
            O => \N__12564\,
            I => \N__12556\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12561\,
            I => \N__12556\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__12556\,
            I => \N__12553\
        );

    \I__2177\ : Sp12to4
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__2176\ : Odrv12
    port map (
            O => \N__12550\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__12538\,
            I => \Lab_UT.dictrl.G_25_i_o3_4\
        );

    \I__2171\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12532\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12532\,
            I => \Lab_UT.dictrl.G_25_i_o3_5\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12529\,
            I => \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__12526\,
            I => \Lab_UT.dictrl.N_11_cascade_\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12512\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12519\,
            I => \N__12512\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12518\,
            I => \N__12507\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12507\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12512\,
            I => \N__12504\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12507\,
            I => \N__12501\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__12504\,
            I => \N__12496\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__12501\,
            I => \N__12496\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__12496\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__12493\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12490\,
            I => \N__12486\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12483\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12486\,
            I => \N__12479\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12483\,
            I => \N__12476\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12473\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__12479\,
            I => \N__12470\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__12476\,
            I => \N__12465\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12465\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__12470\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__12465\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__12460\,
            I => \N__12453\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12450\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12447\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12442\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12442\
        );

    \I__2141\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12439\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__12450\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__12447\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12442\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12439\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12427\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__12427\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__12424\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12418\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12418\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12412\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12412\,
            I => \N__12409\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__12409\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__12406\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12400\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12400\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12384\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12384\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12394\,
            I => \N__12384\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12391\,
            I => \N__12379\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12384\,
            I => \N__12379\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__12379\,
            I => \N__12376\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__12376\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12370\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__12370\,
            I => \N__12365\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12362\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12359\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__12365\,
            I => \N__12354\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12362\,
            I => \N__12354\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12359\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__12354\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12346\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12346\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__12343\,
            I => \Lab_UT.didp.countrce4.q_5_0_cascade_\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12336\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__12336\,
            I => \N__12330\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12327\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__12330\,
            I => \N__12324\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12327\,
            I => \N__12321\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__12324\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__12321\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2098\ : CEMux
    port map (
            O => \N__12316\,
            I => \N__12313\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12310\
        );

    \I__2096\ : Span4Mux_v
    port map (
            O => \N__12310\,
            I => \N__12307\
        );

    \I__2095\ : Span4Mux_h
    port map (
            O => \N__12307\,
            I => \N__12304\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__12304\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__12301\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_\
        );

    \I__2092\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12295\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__12295\,
            I => \N__12292\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__12292\,
            I => \Lab_UT.didp.countrce2.N_96\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__12289\,
            I => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_\
        );

    \I__2088\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12282\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12278\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12282\,
            I => \N__12275\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12272\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12269\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__12275\,
            I => \N__12266\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__12269\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__12266\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__12263\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \N__12249\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__12255\,
            I => \N__12245\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12234\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12234\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12234\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12234\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12234\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12231\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12234\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__12231\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12221\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12218\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12215\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12212\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12218\,
            I => \N__12209\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12206\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12203\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__12209\,
            I => \N__12200\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__12206\,
            I => \N__12197\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__12203\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__12200\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__12197\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12187\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12184\
        );

    \I__2054\ : Span4Mux_h
    port map (
            O => \N__12184\,
            I => \N__12181\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__12181\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12175\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12175\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12169\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12163\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12163\,
            I => \N__12160\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__12160\,
            I => \N__12157\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__12157\,
            I => \uu2.N_149\
        );

    \I__2044\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12151\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12151\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12148\,
            I => \N__12145\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12142\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12142\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12139\,
            I => \N__12136\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12136\,
            I => \uu2.N_25\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__12133\,
            I => \N__12130\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12124\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12124\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__12124\,
            I => \N__12118\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12111\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12111\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12111\
        );

    \I__2030\ : Odrv12
    port map (
            O => \N__12118\,
            I => \Lab_UT.didp.un24_ce_3\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12111\,
            I => \Lab_UT.didp.un24_ce_3\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__12106\,
            I => \N__12098\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12091\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12080\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12080\
        );

    \I__2023\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12080\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12080\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12080\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__12094\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12091\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12080\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12070\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12070\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__12067\,
            I => \N__12064\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12061\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__12061\,
            I => \N__12058\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__12058\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12052\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12052\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__12049\,
            I => \N__12046\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12043\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__12043\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__12040\,
            I => \uu2.N_24_cascade_\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12031\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12031\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12031\,
            I => \uu2.N_31_i\
        );

    \I__2002\ : InMux
    port map (
            O => \N__12028\,
            I => \N__12025\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12025\,
            I => \uu2.N_166\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__12022\,
            I => \uu2.bitmap_pmux_27_ns_1_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12016\,
            I => \uu2.N_26\
        );

    \I__1997\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12010\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__12007\
        );

    \I__1995\ : Span4Mux_s2_v
    port map (
            O => \N__12007\,
            I => \N__12004\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__12004\,
            I => \uu2.N_404\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12001\,
            I => \N__11998\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11998\,
            I => \N__11995\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__11995\,
            I => \N__11992\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__11992\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11978\
        );

    \I__1987\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11978\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11975\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__11983\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11978\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__11975\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11965\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__11965\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__11962\,
            I => \uu2.N_14_cascade_\
        );

    \I__1979\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11956\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__11956\,
            I => \uu2.bitmap_pmux_sn_N_54_mux\
        );

    \I__1977\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11950\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__11950\,
            I => \uu2.bitmap_RNI2Q8F1Z0Z_111\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11940\
        );

    \I__1974\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11933\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11933\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11933\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11930\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__11940\,
            I => \N__11927\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__11933\,
            I => \N__11924\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__11930\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__11927\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__11924\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11914\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11914\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__11911\,
            I => \N__11907\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11902\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11902\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__11902\,
            I => bu_rx_data_fast_5
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__11899\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__11895\,
            I => \N__11887\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__11894\,
            I => \N__11883\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__11893\,
            I => \N__11878\
        );

    \I__1954\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11875\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11862\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11862\
        );

    \I__1951\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11862\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11862\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11862\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11862\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__11875\,
            I => \N__11859\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11856\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__11859\,
            I => \N__11851\
        );

    \I__1944\ : Span4Mux_s0_v
    port map (
            O => \N__11856\,
            I => \N__11851\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__11851\,
            I => \uu2.N_37\
        );

    \I__1942\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__11842\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__11839\,
            I => \resetGen.escKeyZ0Z_4_cascade_\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11821\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11821\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11821\
        );

    \I__1935\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11821\
        );

    \I__1934\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11821\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__11818\,
            I => \N__11815\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__11815\,
            I => \resetGen.escKeyZ0\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11809\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11809\,
            I => \resetGen.escKeyZ0Z_5\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11803\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__11803\,
            I => \Lab_UT.dictrl.g1_0Z0Z_5\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11800\,
            I => \N__11797\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11797\,
            I => \N__11794\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__11794\,
            I => \Lab_UT.dictrl.g1_4_0\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__11791\,
            I => \Lab_UT.dictrl.g1_5_0_cascade_\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__11788\,
            I => \Lab_UT.dictrl.G_25_i_o3_3_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11782\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11782\,
            I => \Lab_UT.dictrl.g0_5_3_0\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11771\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11768\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11765\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11771\,
            I => \Lab_UT.dispString.N_144\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__11768\,
            I => \Lab_UT.dispString.N_144\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__11765\,
            I => \Lab_UT.dispString.N_144\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11755\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__11755\,
            I => \Lab_UT.dispString.N_124\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__11752\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11740\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11737\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11734\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11731\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11740\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11737\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__11734\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__11731\,
            I => \Lab_UT.dispString.N_95\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11719\,
            I => \Lab_UT.dispString.N_102\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__11716\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11710\,
            I => \N__11707\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__11707\,
            I => \N__11704\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__11704\,
            I => \N__11699\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11694\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11694\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11699\,
            I => \L3_tx_data_0\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11694\,
            I => \L3_tx_data_0\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11681\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11681\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11678\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11675\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11681\,
            I => \N__11672\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__11678\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__11675\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__11672\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11661\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \N__11658\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11650\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11647\
        );

    \I__1877\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11642\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11642\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__11655\,
            I => \N__11638\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11634\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__11653\,
            I => \N__11631\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11626\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11647\,
            I => \N__11626\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11623\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11618\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11618\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11611\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11611\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11611\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__11626\,
            I => \N__11608\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__11623\,
            I => \oneSecStrb\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11618\,
            I => \oneSecStrb\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11611\,
            I => \oneSecStrb\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__11608\,
            I => \oneSecStrb\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__11590\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_1\
        );

    \I__1855\ : CEMux
    port map (
            O => \N__11587\,
            I => \N__11584\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11584\,
            I => \N__11581\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__11578\,
            I => \Lab_UT.didp.regrce2.LdAStens_0\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11568\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11574\,
            I => \N__11568\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11562\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__11568\,
            I => \N__11559\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11552\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11552\
        );

    \I__1845\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11552\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11562\,
            I => \N__11549\
        );

    \I__1843\ : Span4Mux_h
    port map (
            O => \N__11559\,
            I => \N__11544\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11552\,
            I => \N__11544\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__11549\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__11544\,
            I => \Lab_UT.dispString.un42_dOutP_1\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \Lab_UT.dispString.N_102_cascade_\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11533\,
            I => \N__11529\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11526\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__11529\,
            I => \G_186\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11526\,
            I => \G_186\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11518\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__11518\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_2\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__11515\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__11509\,
            I => \N__11505\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__11508\,
            I => \N__11501\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__11505\,
            I => \N__11498\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11493\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11493\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__11498\,
            I => \L3_tx_data_2\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11493\,
            I => \L3_tx_data_2\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11484\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11481\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11478\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11481\,
            I => \N__11472\
        );

    \I__1818\ : Span4Mux_s3_v
    port map (
            O => \N__11478\,
            I => \N__11472\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11469\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__11472\,
            I => \L3_tx_data_rdy\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11469\,
            I => \L3_tx_data_rdy\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11456\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11453\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11450\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__11456\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__11453\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11450\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11435\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11432\
        );

    \I__1804\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11429\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__11435\,
            I => \uu2.un1_w_user_crZ0Z_3\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__11432\,
            I => \uu2.un1_w_user_crZ0Z_3\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__11429\,
            I => \uu2.un1_w_user_crZ0Z_3\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11419\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__11416\,
            I => \N__11404\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11401\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11398\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11395\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11392\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11387\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11387\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11380\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11380\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11380\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__11404\,
            I => \G_179\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11401\,
            I => \G_179\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__11398\,
            I => \G_179\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11395\,
            I => \G_179\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__11392\,
            I => \G_179\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11387\,
            I => \G_179\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11380\,
            I => \G_179\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11359\,
            I => \N__11355\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \N__11349\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__11355\,
            I => \N__11340\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11335\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11335\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11332\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11325\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11325\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11325\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11316\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11316\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11316\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11343\,
            I => \N__11316\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__11340\,
            I => \G_181\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11335\,
            I => \G_181\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11332\,
            I => \G_181\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11325\,
            I => \G_181\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__11316\,
            I => \G_181\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11305\,
            I => \N__11302\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11302\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__11299\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__11290\,
            I => \Lab_UT.didp.countrce1.q_5_3\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__1752\ : Span4Mux_v
    port map (
            O => \N__11278\,
            I => \N__11275\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__11275\,
            I => \Lab_UT.dispString.N_137\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11269\,
            I => \N__11265\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11262\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__11265\,
            I => \uu0_sec_clkD\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11262\,
            I => \uu0_sec_clkD\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__11257\,
            I => \Lab_UT.dispString.N_143_cascade_\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11247\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11244\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11247\,
            I => \N__11239\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11239\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__11236\,
            I => \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11230\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11226\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11223\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__11226\,
            I => \N__11220\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11217\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__11220\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__1731\ : Odrv12
    port map (
            O => \N__11217\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11212\,
            I => \N__11209\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11209\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11200\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11197\
        );

    \I__1725\ : Sp12to4
    port map (
            O => \N__11197\,
            I => \N__11194\
        );

    \I__1724\ : Span12Mux_s3_v
    port map (
            O => \N__11194\,
            I => \N__11189\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11184\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11184\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__11189\,
            I => \Lab_UT.didp.ce_12_1\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11184\,
            I => \Lab_UT.didp.ce_12_1\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \Lab_UT.didp.ce_12_1_cascade_\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__11176\,
            I => \Lab_UT.didp.ce_12_3_cascade_\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11161\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11161\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11161\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11161\,
            I => \Lab_UT.didp.countrce1.ce_12_1_1\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__11155\,
            I => \Lab_UT.didp.countrce3.un13_qPone_cascade_\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__11152\,
            I => \Lab_UT.didp.countrce3.q_5_2_cascade_\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11145\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11142\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11145\,
            I => \N__11139\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11136\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__11139\,
            I => \N__11132\
        );

    \I__1704\ : Span4Mux_s2_v
    port map (
            O => \N__11136\,
            I => \N__11125\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \N__11121\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__11132\,
            I => \N__11116\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11113\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__11130\,
            I => \N__11107\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__11129\,
            I => \N__11104\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11101\
        );

    \I__1697\ : Sp12to4
    port map (
            O => \N__11125\,
            I => \N__11098\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11089\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11089\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11089\
        );

    \I__1693\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11089\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__11116\,
            I => \N__11084\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11084\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11073\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11073\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11073\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11073\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11073\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11070\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__11098\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11089\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__11084\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11073\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11070\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11056\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11056\,
            I => \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__11053\,
            I => \N__11050\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11044\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11044\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11044\,
            I => \N__11041\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__11041\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__11038\,
            I => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\
        );

    \I__1671\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11032\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__11032\,
            I => \uu2.bitmap_pmux_sn_i5_mux\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11025\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11022\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11025\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__11022\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__11017\,
            I => \uu2.bitmap_pmux_sn_N_15_cascade_\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11011\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__11011\,
            I => \uu2.N_401\
        );

    \I__1662\ : InMux
    port map (
            O => \N__11008\,
            I => \N__11005\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11005\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10984\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10984\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10984\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10984\
        );

    \I__1656\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10984\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10984\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__10984\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10974\
        );

    \I__1651\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10971\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10974\,
            I => \G_182\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__10971\,
            I => \G_182\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10957\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10957\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10957\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__10957\,
            I => \G_183\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__10954\,
            I => \G_182_cascade_\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10948\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10948\,
            I => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__10945\,
            I => \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10937\
        );

    \I__1639\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10932\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10932\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__10937\,
            I => \Lab_UT.dictrl.alarmstateZ0Z8\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__10932\,
            I => \Lab_UT.dictrl.alarmstateZ0Z8\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__10927\,
            I => \Lab_UT.dictrl.g1_0_4_0_cascade_\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10921\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__10921\,
            I => \Lab_UT.dictrl.g1_0Z0Z_1\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__10918\,
            I => \Lab_UT.dictrl.g0_5_4_0_cascade_\
        );

    \I__1631\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10911\
        );

    \I__1630\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10908\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__10911\,
            I => \G_188\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__10908\,
            I => \G_188\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10900\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__10900\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_3\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__10897\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10891\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__10891\,
            I => \N__10888\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__10888\,
            I => \N__10883\
        );

    \I__1621\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10878\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10878\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__10883\,
            I => \L3_tx_data_3\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10878\,
            I => \L3_tx_data_3\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__10873\,
            I => \G_186_cascade_\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10864\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10864\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__10864\,
            I => \G_187\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__10861\,
            I => \G_187_cascade_\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10855\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__10855\,
            I => \Lab_UT.dispString.dOutP_1_iv_i_1_4\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__10852\,
            I => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\
        );

    \I__1609\ : IoInMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10842\
        );

    \I__1607\ : SRMux
    port map (
            O => \N__10845\,
            I => \N__10839\
        );

    \I__1606\ : IoSpan4Mux
    port map (
            O => \N__10842\,
            I => \N__10835\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10832\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__10838\,
            I => \N__10829\
        );

    \I__1603\ : Span4Mux_s1_v
    port map (
            O => \N__10835\,
            I => \N__10824\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__10832\,
            I => \N__10824\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10821\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__10824\,
            I => \N__10816\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10821\,
            I => \N__10813\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10810\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10807\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__10816\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1595\ : Odrv12
    port map (
            O => \N__10813\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10810\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10807\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__10798\,
            I => \uu2.un1_w_user_lfZ0Z_4_cascade_\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10789\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10789\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10786\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__10786\,
            I => \uu2.un20_w_addr_userZ0Z_1\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10780\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__1585\ : Span12Mux_s3_v
    port map (
            O => \N__10777\,
            I => \N__10772\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10767\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10767\
        );

    \I__1582\ : Odrv12
    port map (
            O => \N__10772\,
            I => \L3_tx_data_1\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10767\,
            I => \L3_tx_data_1\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10759\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10756\
        );

    \I__1578\ : Span4Mux_s3_v
    port map (
            O => \N__10756\,
            I => \N__10751\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10755\,
            I => \N__10746\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10746\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__10751\,
            I => \L3_tx_data_4\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10746\,
            I => \L3_tx_data_4\
        );

    \I__1573\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10737\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__10740\,
            I => \N__10734\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10730\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10727\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10724\
        );

    \I__1568\ : Odrv12
    port map (
            O => \N__10730\,
            I => \L3_tx_data_6\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10727\,
            I => \L3_tx_data_6\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__10724\,
            I => \L3_tx_data_6\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10714\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__10714\,
            I => \uu2.un1_w_user_lfZ0Z_3\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__10711\,
            I => \N__10708\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10705\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10705\,
            I => \N__10702\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__10702\,
            I => \Lab_UT.dispString.N_140\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10695\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__10689\,
            I => \N__10682\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10679\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10676\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__10682\,
            I => \L3_tx_data_5\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__10679\,
            I => \L3_tx_data_5\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10676\,
            I => \L3_tx_data_5\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__10669\,
            I => \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10662\
        );

    \I__1547\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10659\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__10662\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10659\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10651\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10651\,
            I => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10645\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10645\,
            I => \uu2.w_addr_displaying_RNI0NG56Z0Z_4\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10639\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10639\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10632\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10629\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10632\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10629\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10621\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10621\,
            I => \N__10618\
        );

    \I__1532\ : Sp12to4
    port map (
            O => \N__10618\,
            I => \N__10615\
        );

    \I__1531\ : Span12Mux_s10_v
    port map (
            O => \N__10615\,
            I => \N__10612\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__10612\,
            I => \uart_RXD\
        );

    \I__1529\ : SRMux
    port map (
            O => \N__10609\,
            I => \N__10605\
        );

    \I__1528\ : CEMux
    port map (
            O => \N__10608\,
            I => \N__10602\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10605\,
            I => \N__10599\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10602\,
            I => \N__10596\
        );

    \I__1525\ : Span4Mux_s3_h
    port map (
            O => \N__10599\,
            I => \N__10591\
        );

    \I__1524\ : Span4Mux_s0_v
    port map (
            O => \N__10596\,
            I => \N__10591\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__10591\,
            I => \N__10588\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__10588\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10582\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10582\,
            I => \uu2.w_addr_displaying_RNI03P31Z0Z_4\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10579\,
            I => \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10573\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10573\,
            I => \uu2.bitmap_pmux_sn_i7_mux_0\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \uu2.N_406_cascade_\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10561\
        );

    \I__1514\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10561\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10561\,
            I => \uu2.bitmap_pmux\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__10558\,
            I => \uu2.N_383_cascade_\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10555\,
            I => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10549\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10549\,
            I => \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10543\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__10543\,
            I => \uu2.bitmap_pmux_u_1\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__10540\,
            I => \uu2.un28_w_addr_user_i_cascade_\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__10537\,
            I => \N__10533\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__10536\,
            I => \N__10530\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10524\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10524\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10521\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10524\,
            I => \uu2.un51_w_data_displaying_i_a2_1\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10521\,
            I => \uu2.un51_w_data_displaying_i_a2_1\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__10516\,
            I => \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10507\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__10507\,
            I => \uu2.w_data_displaying_2_i_a2_i_a3_2_0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__10504\,
            I => \G_179_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10495\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10488\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10488\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10488\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10495\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10488\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__10483\,
            I => \Lab_UT.un1_idle_5_0_iclkZ0_cascade_\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10476\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10473\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10476\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10473\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10464\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10461\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10464\,
            I => \G_185\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10461\,
            I => \G_185\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10453\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10450\
        );

    \I__1476\ : Span4Mux_h
    port map (
            O => \N__10450\,
            I => \N__10447\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__10447\,
            I => vbuf_tx_data_6
        );

    \I__1474\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10441\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10441\,
            I => \N__10438\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__10438\,
            I => \N__10435\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__10435\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10429\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__10429\,
            I => \N__10426\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__10426\,
            I => vbuf_tx_data_7
        );

    \I__1467\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10420\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10420\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \N__10414\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10411\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10408\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__10408\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__1461\ : CEMux
    port map (
            O => \N__10405\,
            I => \N__10402\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10402\,
            I => \N__10399\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__10399\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__10396\,
            I => \Lab_UT.un1_idle_1_0_iclkZ0_cascade_\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__10393\,
            I => \Lab_UT.dispString.N_117_cascade_\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10390\,
            I => \G_180_cascade_\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__10387\,
            I => \G_181_cascade_\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10381\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10381\,
            I => \G_180\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__10378\,
            I => \Lab_UT.dictrl.alarmstate_1_0_cascade_\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__10374\,
            I => \N__10366\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10362\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10359\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10356\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10351\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10351\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10348\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10359\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__10356\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__10351\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10348\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10334\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10326\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10326\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10323\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10320\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10315\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10315\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10326\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__10323\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10320\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10315\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10300\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10297\
        );

    \I__1425\ : Odrv12
    port map (
            O => \N__10297\,
            I => \uu2.un284_ci\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__10294\,
            I => \Lab_UT.didp.countrce1.q_5_0_cascade_\
        );

    \I__1423\ : CEMux
    port map (
            O => \N__10291\,
            I => \N__10287\
        );

    \I__1422\ : CEMux
    port map (
            O => \N__10290\,
            I => \N__10284\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10287\,
            I => \N__10281\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10284\,
            I => \N__10278\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__10281\,
            I => \N__10275\
        );

    \I__1418\ : Odrv12
    port map (
            O => \N__10278\,
            I => \Lab_UT.didp.regrce3.LdAMones_0\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__10275\,
            I => \Lab_UT.didp.regrce3.LdAMones_0\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10267\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10267\,
            I => \G_184\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__10264\,
            I => \G_184_cascade_\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10261\,
            I => \N__10256\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10248\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10248\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10245\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10238\
        );

    \I__1408\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10238\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10238\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10248\,
            I => \N__10235\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10245\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10238\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__10235\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1402\ : CEMux
    port map (
            O => \N__10228\,
            I => \N__10225\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10222\
        );

    \I__1400\ : Odrv12
    port map (
            O => \N__10222\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10216\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10216\,
            I => \N__10213\
        );

    \I__1397\ : Span4Mux_s0_v
    port map (
            O => \N__10213\,
            I => \N__10210\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__10210\,
            I => \uu2.mem0.w_data_2\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__10207\,
            I => \N__10201\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10198\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10192\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10192\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10189\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10198\,
            I => \N__10186\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10183\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10180\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10189\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__10186\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__10183\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__10180\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__10171\,
            I => \N__10168\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10159\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10156\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10153\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10162\,
            I => \N__10146\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10159\,
            I => \N__10146\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__10156\,
            I => \N__10146\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10153\,
            I => \uu2.un404_ci_0\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__10146\,
            I => \uu2.un404_ci_0\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10133\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10122\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10122\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10122\
        );

    \I__1369\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10122\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10122\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__10133\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10122\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10113\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10104\
        );

    \I__1361\ : Span4Mux_s0_v
    port map (
            O => \N__10107\,
            I => \N__10097\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10097\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10094\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \N__10091\
        );

    \I__1357\ : Span4Mux_v
    port map (
            O => \N__10097\,
            I => \N__10086\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10094\,
            I => \N__10086\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10083\
        );

    \I__1354\ : Span4Mux_s0_v
    port map (
            O => \N__10086\,
            I => \N__10080\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__10083\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__10080\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10072\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10065\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10056\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10056\
        );

    \I__1347\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10056\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10056\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__10065\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__10056\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10045\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10041\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10038\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__10041\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__10038\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10030\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10030\,
            I => \N__10027\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__10027\,
            I => \N__10020\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10011\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10011\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10011\
        );

    \I__1331\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10011\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__10020\,
            I => \uu2.un306_ci\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__10011\,
            I => \uu2.un306_ci\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10006\,
            I => \N__10002\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9998\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9995\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9992\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__1323\ : Span4Mux_s3_h
    port map (
            O => \N__9995\,
            I => \N__9986\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9992\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__9989\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__9986\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__9976\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__9970\,
            I => \uu2.N_34\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__9967\,
            I => \uu2.N_34_cascade_\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9961\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__9961\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9955\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__9955\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9952\,
            I => \N__9949\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9949\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9940\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__9940\,
            I => \uu2.N_31\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \uu2.N_31_cascade_\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__9931\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__9928\,
            I => \N__9923\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9927\,
            I => \N__9917\
        );

    \I__1300\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9917\
        );

    \I__1299\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9914\
        );

    \I__1298\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9911\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9917\,
            I => \N__9908\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__9914\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__9911\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__9908\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__9901\,
            I => \N__9897\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__9900\,
            I => \N__9892\
        );

    \I__1291\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9888\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9883\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9883\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9878\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9878\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9873\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__9883\,
            I => \N__9873\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__9878\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__9873\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__9868\,
            I => \uu2.vbuf_raddr.un448_ci_0_cascade_\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__9865\,
            I => \N__9862\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9858\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9855\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9858\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9855\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9847\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9842\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9837\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9837\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9842\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9837\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__9832\,
            I => \N__9827\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__9831\,
            I => \N__9824\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__9830\,
            I => \N__9821\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9818\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9813\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9813\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9818\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__9813\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__9808\,
            I => \uu2.un404_ci_0_cascade_\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__9805\,
            I => \N__9802\
        );

    \I__1260\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9796\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9789\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9789\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9799\,
            I => \N__9789\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__9796\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__9789\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9778\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__9778\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9772\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__9772\,
            I => \uu2.mem0.w_data_6\
        );

    \I__1249\ : CEMux
    port map (
            O => \N__9769\,
            I => \N__9763\
        );

    \I__1248\ : CEMux
    port map (
            O => \N__9768\,
            I => \N__9760\
        );

    \I__1247\ : CEMux
    port map (
            O => \N__9767\,
            I => \N__9757\
        );

    \I__1246\ : CEMux
    port map (
            O => \N__9766\,
            I => \N__9754\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9763\,
            I => \N__9749\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9760\,
            I => \N__9749\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9746\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9743\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__9749\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1240\ : Odrv12
    port map (
            O => \N__9746\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__9743\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9731\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9726\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9726\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9731\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__9726\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9717\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__9720\,
            I => \N__9713\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9709\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9702\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9702\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9702\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9709\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9702\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1225\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9692\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9687\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9687\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9692\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9687\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9679\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9676\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9669\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9666\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9669\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__9666\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9661\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9653\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9648\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9648\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9653\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__9648\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__1206\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9637\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9634\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__9631\,
            I => \N__9625\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9622\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9615\
        );

    \I__1200\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9615\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9615\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9622\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__9615\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9610\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__9607\,
            I => \N__9603\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__9606\,
            I => \N__9600\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9597\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9597\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9594\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9582\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9582\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9579\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9582\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__9579\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__9574\,
            I => \N__9571\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9561\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9561\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9561\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9558\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__9561\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9558\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__9553\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9546\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9543\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9546\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9543\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__9538\,
            I => \N__9531\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9521\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9521\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9521\
        );

    \I__1168\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9521\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9531\,
            I => \N__9516\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9516\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9521\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__9516\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9505\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9505\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9502\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__9502\,
            I => \resetGen.un241_ci\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__9499\,
            I => \N__9496\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9489\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9489\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9486\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9489\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9486\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__9481\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__9472\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__9469\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__9466\,
            I => \N__9462\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9465\,
            I => \N__9458\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9455\
        );

    \I__1145\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9450\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9445\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9445\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9440\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9440\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9450\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__9445\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__9440\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1137\ : IoInMux
    port map (
            O => \N__9433\,
            I => \N__9430\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__9430\,
            I => \N__9427\
        );

    \I__1135\ : Span12Mux_s4_v
    port map (
            O => \N__9427\,
            I => \N__9424\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__9424\,
            I => \buart.Z_rx.sample\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__9421\,
            I => \N__9418\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9415\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9415\,
            I => \N__9412\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__9412\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9402\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9396\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__9402\,
            I => \N__9393\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9386\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9386\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9386\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__9396\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__9393\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9386\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9374\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9368\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9368\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9374\,
            I => \N__9365\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9362\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9368\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__9365\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9362\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9352\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9352\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9345\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9342\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9345\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__9342\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9333\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9327\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9333\,
            I => \N__9317\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9310\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9310\
        );

    \I__1100\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9310\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9327\,
            I => \N__9307\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9299\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9299\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9299\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9296\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9293\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9290\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9287\
        );

    \I__1091\ : Span4Mux_v
    port map (
            O => \N__9317\,
            I => \N__9284\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9279\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__9307\,
            I => \N__9279\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9276\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__9299\,
            I => \uu0.un4_l_count_0\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9296\,
            I => \uu0.un4_l_count_0\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__9293\,
            I => \uu0.un4_l_count_0\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9290\,
            I => \uu0.un4_l_count_0\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9287\,
            I => \uu0.un4_l_count_0\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__9284\,
            I => \uu0.un4_l_count_0\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__9279\,
            I => \uu0.un4_l_count_0\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__9276\,
            I => \uu0.un4_l_count_0\
        );

    \I__1079\ : IoInMux
    port map (
            O => \N__9259\,
            I => \N__9256\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9256\,
            I => \N__9253\
        );

    \I__1077\ : Span4Mux_s1_h
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__9250\,
            I => \uu0.un11_l_count_i\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9247\,
            I => \N__9244\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__1072\ : Span12Mux_s9_v
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__1071\ : Odrv12
    port map (
            O => \N__9235\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__9229\,
            I => \resetGen.reset_count_2_0_4\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9220\,
            I => \uu0.un99_ci_0\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9212\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9207\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9207\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9212\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9207\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9199\,
            I => \uu0.un44_ci\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__9196\,
            I => \uu0.un44_ci_cascade_\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9188\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9183\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9183\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9188\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9183\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9172\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9161\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9161\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9158\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__9166\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9161\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9158\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__9151\,
            I => \N__9144\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__9150\,
            I => \N__9141\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9132\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9132\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9132\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9132\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9129\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9132\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9129\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__1034\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9114\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9114\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9114\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9111\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__9114\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9111\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__9106\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9092\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9092\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9089\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9086\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9083\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__9089\,
            I => \uu0.un66_ci\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__9086\,
            I => \uu0.un66_ci\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__9083\,
            I => \uu0.un66_ci\
        );

    \I__1018\ : CEMux
    port map (
            O => \N__9076\,
            I => \N__9064\
        );

    \I__1017\ : CEMux
    port map (
            O => \N__9075\,
            I => \N__9064\
        );

    \I__1016\ : CEMux
    port map (
            O => \N__9074\,
            I => \N__9064\
        );

    \I__1015\ : CEMux
    port map (
            O => \N__9073\,
            I => \N__9064\
        );

    \I__1014\ : GlobalMux
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__1013\ : gio2CtrlBuf
    port map (
            O => \N__9061\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9045\
        );

    \I__1010\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9045\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9045\
        );

    \I__1008\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9042\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__9045\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9042\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9030\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9030\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9027\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9030\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9027\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__9022\,
            I => \N__9017\
        );

    \I__999\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9010\
        );

    \I__998\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9010\
        );

    \I__997\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9010\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__9007\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__9007\,
            I => \uu0.un88_ci_3\
        );

    \I__994\ : InMux
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8998\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__8998\,
            I => \uu0.un187_ci_1\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__8995\,
            I => \N__8991\
        );

    \I__990\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8988\
        );

    \I__989\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8981\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8978\
        );

    \I__986\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8975\
        );

    \I__985\ : Span4Mux_s1_h
    port map (
            O => \N__8981\,
            I => \N__8972\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__8978\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__8975\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__8972\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__981\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8962\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8962\,
            I => \uu0.un4_l_count_12\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__8959\,
            I => \N__8954\
        );

    \I__978\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8949\
        );

    \I__977\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8949\
        );

    \I__976\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8946\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__8949\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__8946\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8936\
        );

    \I__972\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8929\
        );

    \I__971\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8929\
        );

    \I__970\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8929\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8926\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__8926\,
            I => \uu0.un198_ci_2\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__8923\,
            I => \N__8920\
        );

    \I__966\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__965\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8909\
        );

    \I__964\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8909\
        );

    \I__963\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8906\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__8914\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__8909\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8906\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__8899\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8892\
        );

    \I__957\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8889\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8892\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__8889\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__8883\,
            I => \N__8873\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__8882\,
            I => \N__8870\
        );

    \I__951\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8863\
        );

    \I__950\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8856\
        );

    \I__949\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8856\
        );

    \I__948\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8856\
        );

    \I__947\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8847\
        );

    \I__946\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8847\
        );

    \I__945\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8847\
        );

    \I__944\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8847\
        );

    \I__943\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8842\
        );

    \I__942\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8842\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8835\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8856\,
            I => \N__8835\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8847\,
            I => \N__8835\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8842\,
            I => \uu0.un110_ci\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__8835\,
            I => \uu0.un110_ci\
        );

    \I__936\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8822\
        );

    \I__935\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8811\
        );

    \I__934\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8811\
        );

    \I__933\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8811\
        );

    \I__932\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8811\
        );

    \I__931\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8811\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8822\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8811\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__928\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8799\
        );

    \I__927\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8794\
        );

    \I__926\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8794\
        );

    \I__925\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8789\
        );

    \I__924\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8789\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__8799\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8794\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__8789\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__8782\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__919\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8770\
        );

    \I__918\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8770\
        );

    \I__917\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8770\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__8770\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__915\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8760\
        );

    \I__914\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8751\
        );

    \I__913\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8751\
        );

    \I__912\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8751\
        );

    \I__911\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8751\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8746\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8746\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__8746\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__907\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8737\
        );

    \I__906\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8734\
        );

    \I__905\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8729\
        );

    \I__904\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8729\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8737\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8734\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8729\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__8722\,
            I => \uu0.un165_ci_0_cascade_\
        );

    \I__899\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8713\
        );

    \I__898\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8713\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8713\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__8710\,
            I => \N__8707\
        );

    \I__895\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8701\
        );

    \I__894\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8698\
        );

    \I__893\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8695\
        );

    \I__892\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8692\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__8701\,
            I => \N__8689\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8698\,
            I => \uu0.un154_ci_9\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__8695\,
            I => \uu0.un154_ci_9\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8692\,
            I => \uu0.un154_ci_9\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__8689\,
            I => \uu0.un154_ci_9\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__8680\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__885\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8668\
        );

    \I__884\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8668\
        );

    \I__883\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8668\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__8668\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__881\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8659\
        );

    \I__880\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8652\
        );

    \I__879\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8652\
        );

    \I__878\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8652\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__8659\,
            I => \N__8649\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__8652\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__8649\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__8644\,
            I => \N__8639\
        );

    \I__873\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8636\
        );

    \I__872\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8631\
        );

    \I__871\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8631\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8636\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8631\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \N__8620\
        );

    \I__867\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8608\
        );

    \I__866\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8608\
        );

    \I__865\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8608\
        );

    \I__864\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8608\
        );

    \I__863\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8608\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8608\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__861\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8598\
        );

    \I__860\ : InMux
    port map (
            O => \N__8604\,
            I => \N__8598\
        );

    \I__859\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8595\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8598\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8595\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__8590\,
            I => \N__8585\
        );

    \I__855\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8582\
        );

    \I__854\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8579\
        );

    \I__853\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8576\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8582\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8579\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8576\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__8569\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__848\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8563\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8563\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__846\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8554\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__8559\,
            I => \N__8551\
        );

    \I__844\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8548\
        );

    \I__843\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8545\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8542\
        );

    \I__841\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8539\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8548\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__8545\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__8542\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8539\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__836\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8527\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__834\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8521\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__8521\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__832\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8513\
        );

    \I__831\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8508\
        );

    \I__830\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8508\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8513\,
            I => \N__8505\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8508\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__8505\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__826\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8497\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__8497\,
            I => vbuf_tx_data_2
        );

    \I__824\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8491\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8491\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__822\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8485\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8485\,
            I => vbuf_tx_data_3
        );

    \I__820\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8479\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__818\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8473\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8473\,
            I => vbuf_tx_data_4
        );

    \I__816\ : InMux
    port map (
            O => \N__8470\,
            I => \N__8467\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8467\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__814\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8461\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8461\,
            I => vbuf_tx_data_5
        );

    \I__812\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8455\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8455\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__8452\,
            I => \uu2.vbuf_count.un328_ci_3_cascade_\
        );

    \I__809\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8446\,
            I => \uu2.un350_ci\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__8443\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__806\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8437\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8437\,
            I => \uu2.r_data_wire_3\
        );

    \I__804\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8431\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8431\,
            I => \uu2.r_data_wire_4\
        );

    \I__802\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8425\,
            I => \uu2.r_data_wire_5\
        );

    \I__800\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8419\,
            I => \uu2.r_data_wire_6\
        );

    \I__798\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8413\,
            I => \uu2.r_data_wire_7\
        );

    \I__796\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8407\,
            I => vbuf_tx_data_0
        );

    \I__794\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8401\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__792\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8395\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8395\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__790\ : IoInMux
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__788\ : Span12Mux_s1_h
    port map (
            O => \N__8386\,
            I => \N__8383\
        );

    \I__787\ : Odrv12
    port map (
            O => \N__8383\,
            I => o_serial_data_c
        );

    \I__786\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8377\,
            I => vbuf_tx_data_1
        );

    \I__784\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8371\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__782\ : InMux
    port map (
            O => \N__8368\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__781\ : InMux
    port map (
            O => \N__8365\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__8362\,
            I => \N__8357\
        );

    \I__779\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8352\
        );

    \I__778\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8343\
        );

    \I__777\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8343\
        );

    \I__776\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8343\
        );

    \I__775\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8343\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8352\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8343\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__772\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8335\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__770\ : InMux
    port map (
            O => \N__8332\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__769\ : InMux
    port map (
            O => \N__8329\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__767\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__766\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8310\
        );

    \I__765\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8310\
        );

    \I__764\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8310\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8317\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8310\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__760\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8299\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__758\ : InMux
    port map (
            O => \N__8296\,
            I => \N__8285\
        );

    \I__757\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8285\
        );

    \I__756\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8285\
        );

    \I__755\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8282\
        );

    \I__754\ : InMux
    port map (
            O => \N__8292\,
            I => \N__8279\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8276\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__8282\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8279\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__8276\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__749\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8266\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8266\,
            I => \uu2.r_data_wire_0\
        );

    \I__747\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8260\,
            I => \uu2.r_data_wire_1\
        );

    \I__745\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8254\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__8254\,
            I => \uu2.r_data_wire_2\
        );

    \I__743\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8244\
        );

    \I__742\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8237\
        );

    \I__741\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8237\
        );

    \I__740\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8237\
        );

    \I__739\ : InMux
    port map (
            O => \N__8247\,
            I => \N__8233\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8244\,
            I => \N__8228\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8237\,
            I => \N__8228\
        );

    \I__736\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8225\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8233\,
            I => \N__8222\
        );

    \I__734\ : Odrv12
    port map (
            O => \N__8228\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8225\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__8222\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__731\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8208\
        );

    \I__730\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8199\
        );

    \I__729\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8199\
        );

    \I__728\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8199\
        );

    \I__727\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8199\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8208\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__8199\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__8194\,
            I => \buart.Z_rx.idle_0_cascade_\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__8191\,
            I => \buart.Z_rx.valid_0_cascade_\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__8188\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__8185\,
            I => \buart.Z_rx.N_27_0_i_cascade_\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__8182\,
            I => \uu0.un143_ci_0_cascade_\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__8179\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__718\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8173\,
            I => \uu0.un4_l_count_18\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__8170\,
            I => \uu0.un4_l_count_16_cascade_\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__8167\,
            I => \N__8162\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__8166\,
            I => \N__8159\
        );

    \I__713\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8152\
        );

    \I__712\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8152\
        );

    \I__711\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8152\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__8152\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__708\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8134\
        );

    \I__707\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8134\
        );

    \I__706\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8134\
        );

    \I__705\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8134\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__8134\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__8131\,
            I => \N__8127\
        );

    \I__702\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8121\
        );

    \I__701\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8121\
        );

    \I__700\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8118\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__8121\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__8118\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__697\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8110\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8110\,
            I => \uu0.un4_l_count_13\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__8107\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__8104\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__693\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8089\
        );

    \I__692\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8089\
        );

    \I__691\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8089\
        );

    \I__690\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8089\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__8089\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__688\ : IoInMux
    port map (
            O => \N__8086\,
            I => \N__8083\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__8083\,
            I => \N__8080\
        );

    \I__686\ : Span12Mux_s9_v
    port map (
            O => \N__8080\,
            I => \N__8077\
        );

    \I__685\ : Odrv12
    port map (
            O => \N__8077\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__684\ : IoInMux
    port map (
            O => \N__8074\,
            I => \N__8071\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__682\ : IoSpan4Mux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__8065\,
            I => clk_in_c
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__22339\
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__22342\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__22346\
        );

    \INVuu2.bitmap_215C\ : INV
    port map (
            O => \INVuu2.bitmap_215C_net\,
            I => \N__22321\
        );

    \INVuu2.w_addr_displaying_7C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_7C_net\,
            I => \N__22338\
        );

    \INVuu2.w_addr_displaying_ness_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_ness_6C_net\,
            I => \N__22341\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__22320\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__22325\
        );

    \INVuu2.bitmap_40C\ : INV
    port map (
            O => \INVuu2.bitmap_40C_net\,
            I => \N__22332\
        );

    \INVuu2.w_addr_displaying_fast_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_8C_net\,
            I => \N__22337\
        );

    \INVuu2.bitmap_197C\ : INV
    port map (
            O => \INVuu2.bitmap_197C_net\,
            I => \N__22315\
        );

    \INVuu2.w_addr_displaying_1_rep1_nesrC\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            I => \N__22323\
        );

    \INVuu2.w_addr_user_2C\ : INV
    port map (
            O => \INVuu2.w_addr_user_2C_net\,
            I => \N__22327\
        );

    \INVuu2.w_addr_displaying_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_3C_net\,
            I => \N__22331\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__22348\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8086\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9433\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9259\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12723\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.l_count_8_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8588\,
            in2 => \_gnd_net_\,
            in3 => \N__8449\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22328\,
            ce => 'H',
            sr => \N__20953\
        );

    \uu2.l_count_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10372\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22328\,
            ce => 'H',
            sr => \N__20953\
        );

    \uu2.l_count_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10337\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22328\,
            ce => 'H',
            sr => \N__20953\
        );

    \uu0.l_precount_0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8236\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22328\,
            ce => 'H',
            sr => \N__20953\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8704\,
            in1 => \N__8557\,
            in2 => \_gnd_net_\,
            in3 => \N__8743\,
            lcout => \uu0.un187_ci_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI04591_10_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8098\,
            in1 => \N__8825\,
            in2 => \N__8559\,
            in3 => \N__9169\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2GS72_4_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8247\,
            in1 => \N__8740\,
            in2 => \N__8107\,
            in3 => \N__9052\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_10_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8101\,
            in1 => \N__8806\,
            in2 => \N__8884\,
            in3 => \N__8828\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => \N__9074\,
            sr => \N__20949\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8826\,
            in1 => \N__8804\,
            in2 => \N__8131\,
            in3 => \N__8099\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8741\,
            in1 => \N__8558\,
            in2 => \N__8104\,
            in3 => \N__8881\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => \N__9074\,
            sr => \N__20949\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8827\,
            in1 => \N__8805\,
            in2 => \_gnd_net_\,
            in3 => \N__8100\,
            lcout => OPEN,
            ltout => \uu0.un143_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_11_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__8877\,
            in1 => \N__8130\,
            in2 => \N__8182\,
            in3 => \N__9323\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => \N__9074\,
            sr => \N__20949\
        );

    \uu0.l_count_8_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8829\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => \N__9074\,
            sr => \N__20949\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8211\,
            in1 => \N__9035\,
            in2 => \N__8166\,
            in3 => \N__9121\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI96A32_18_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8665\,
            in1 => \N__8895\,
            in2 => \N__8179\,
            in3 => \N__8994\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_11_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8113\,
            in1 => \N__8176\,
            in2 => \N__8170\,
            in3 => \N__8965\,
            lcout => \uu0.un4_l_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_2_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__8213\,
            in1 => \N__8145\,
            in2 => \_gnd_net_\,
            in3 => \N__8249\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \N__20951\
        );

    \uu0.l_precount_3_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8250\,
            in1 => \N__8165\,
            in2 => \N__8149\,
            in3 => \N__8214\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \N__20951\
        );

    \uu0.delay_line_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8212\,
            in1 => \N__8144\,
            in2 => \N__8167\,
            in3 => \N__8248\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \N__20951\
        );

    \uu0.l_count_RNI2CNU_11_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8143\,
            in1 => \N__8126\,
            in2 => \N__9150\,
            in3 => \N__8917\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9349\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22300\,
            ce => 'H',
            sr => \N__20952\
        );

    \uu0.l_precount_1_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8251\,
            in2 => \_gnd_net_\,
            in3 => \N__8215\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22300\,
            ce => 'H',
            sr => \N__20952\
        );

    \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8322\,
            in1 => \N__9401\,
            in2 => \N__8362\,
            in3 => \N__8295\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8355\,
            in2 => \_gnd_net_\,
            in3 => \N__8320\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__9399\,
            in2 => \N__8194\,
            in3 => \N__8296\,
            lcout => \buart.Z_rx.idle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8321\,
            in2 => \_gnd_net_\,
            in3 => \N__9453\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8356\,
            in1 => \N__9400\,
            in2 => \N__8191\,
            in3 => \N__8294\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8188\,
            in3 => \N__13784\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => \buart.Z_rx.N_27_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__8360\,
            in1 => \N__8338\,
            in2 => \N__8185\,
            in3 => \N__13759\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22291\,
            ce => \N__9768\,
            sr => \N__20956\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8292\,
            in2 => \_gnd_net_\,
            in3 => \N__8368\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9409\,
            in3 => \N__8365\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8361\,
            in2 => \_gnd_net_\,
            in3 => \N__8332\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__9373\,
            in1 => \N__13757\,
            in2 => \N__8326\,
            in3 => \N__8329\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__9766\,
            sr => \N__20959\
        );

    \buart.Z_rx.bitcount_es_1_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__9379\,
            in1 => \N__8293\,
            in2 => \N__8305\,
            in3 => \N__13760\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22277\,
            ce => \N__9769\,
            sr => \N__20961\
        );

    \uu2.r_data_reg_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8263\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8440\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8434\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8428\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8422\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21708\,
            in1 => \N__8374\,
            in2 => \_gnd_net_\,
            in3 => \N__8410\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_0_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8404\,
            in2 => \_gnd_net_\,
            in3 => \N__21706\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.uart_tx_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8398\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_2_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8494\,
            in1 => \N__21709\,
            in2 => \_gnd_net_\,
            in3 => \N__8380\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_3_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21710\,
            in1 => \N__8482\,
            in2 => \_gnd_net_\,
            in3 => \N__8500\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_4_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8488\,
            in1 => \N__8470\,
            in2 => \_gnd_net_\,
            in3 => \N__21711\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_5_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21712\,
            in1 => \N__8458\,
            in2 => \_gnd_net_\,
            in3 => \N__8476\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \buart.Z_tx.shifter_6_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10444\,
            in1 => \N__21713\,
            in2 => \_gnd_net_\,
            in3 => \N__8464\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => \N__21621\,
            sr => \N__20964\
        );

    \uu0.sec_clk_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13546\,
            in2 => \_gnd_net_\,
            in3 => \N__9336\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22335\,
            ce => 'H',
            sr => \N__20962\
        );

    \uu2.vram_rd_clk_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14347\,
            in2 => \_gnd_net_\,
            in3 => \N__8518\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22335\,
            ce => 'H',
            sr => \N__20962\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8623\,
            in2 => \_gnd_net_\,
            in3 => \N__8604\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => \uu2.vbuf_count.un328_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10005\,
            in1 => \N__10070\,
            in2 => \N__8452\,
            in3 => \N__10023\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__8517\,
            in1 => \N__8643\,
            in2 => \N__8443\,
            in3 => \N__8589\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__20960\
        );

    \uu2.l_count_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8624\,
            in1 => \N__10025\,
            in2 => \_gnd_net_\,
            in3 => \N__8516\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__20960\
        );

    \uu2.l_count_5_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10026\,
            in1 => \N__8625\,
            in2 => \_gnd_net_\,
            in3 => \N__8605\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__20960\
        );

    \uu2.l_count_6_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10044\,
            in1 => \N__10071\,
            in2 => \_gnd_net_\,
            in3 => \N__10024\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__20960\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10068\,
            in1 => \N__8619\,
            in2 => \N__8644\,
            in3 => \N__10331\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_9_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10332\,
            in1 => \N__8642\,
            in2 => \N__8626\,
            in3 => \N__10069\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIFGGK1_3_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8603\,
            in1 => \N__10006\,
            in2 => \N__8590\,
            in3 => \N__8777\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10365\,
            in1 => \N__8763\,
            in2 => \N__8569\,
            in3 => \N__8566\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8984\,
            in1 => \N__8560\,
            in2 => \N__8710\,
            in3 => \N__8742\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8530\,
            in1 => \N__8765\,
            in2 => \N__10374\,
            in3 => \N__8524\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__10306\,
            in1 => \N__8767\,
            in2 => \N__8782\,
            in3 => \N__8779\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \N__20958\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8764\,
            in1 => \N__8778\,
            in2 => \N__10373\,
            in3 => \N__10333\,
            lcout => \uu2.un306_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10305\,
            in2 => \_gnd_net_\,
            in3 => \N__8766\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \N__20958\
        );

    \uu0.l_count_RNIFAQ9_13_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8718\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9020\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8705\,
            in2 => \_gnd_net_\,
            in3 => \N__8676\,
            lcout => OPEN,
            ltout => \uu0.un165_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_13_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8719\,
            in1 => \N__8866\,
            in2 => \N__8722\,
            in3 => \N__9331\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22317\,
            ce => \N__9076\,
            sr => \N__20954\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9099\,
            in1 => \N__8662\,
            in2 => \N__9022\,
            in3 => \N__9217\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_12_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8677\,
            in1 => \N__8706\,
            in2 => \N__8680\,
            in3 => \N__9330\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22317\,
            ce => \N__9076\,
            sr => \N__20954\
        );

    \uu0.l_count_6_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__9021\,
            in1 => \N__9337\,
            in2 => \N__9103\,
            in3 => \N__8664\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22317\,
            ce => \N__9076\,
            sr => \N__20954\
        );

    \uu0.l_count_15_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__9004\,
            in1 => \N__8867\,
            in2 => \N__8995\,
            in3 => \N__9332\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22317\,
            ce => \N__9076\,
            sr => \N__20954\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8802\,
            in1 => \N__9215\,
            in2 => \N__8959\,
            in3 => \N__9191\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__8939\,
            in1 => \N__8869\,
            in2 => \N__8923\,
            in3 => \N__9324\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.l_count_17_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8919\,
            in1 => \N__8940\,
            in2 => \N__8882\,
            in3 => \N__8958\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8957\,
            in1 => \N__8868\,
            in2 => \N__8941\,
            in3 => \N__8918\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9321\,
            in2 => \N__8899\,
            in3 => \N__8896\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.l_count_3_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9192\,
            in1 => \N__9202\,
            in2 => \N__9178\,
            in3 => \N__9326\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.l_count_9_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__8803\,
            in1 => \_gnd_net_\,
            in2 => \N__8883\,
            in3 => \N__8830\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.l_count_7_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9216\,
            in1 => \N__9098\,
            in2 => \N__9226\,
            in3 => \N__9325\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22309\,
            ce => \N__9075\,
            sr => \N__20950\
        );

    \uu0.l_count_0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9322\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => \N__9073\,
            sr => \N__20955\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__9123\,
            in1 => \N__9147\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.un44_ci\,
            ltout => \uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9196\,
            in3 => \N__9171\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => \N__9073\,
            sr => \N__20955\
        );

    \uu0.l_count_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__9124\,
            in1 => \N__9149\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => \N__9073\,
            sr => \N__20955\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9193\,
            in1 => \N__9170\,
            in2 => \N__9151\,
            in3 => \N__9122\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_4_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9320\,
            in2 => \N__9106\,
            in3 => \N__9054\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => \N__9073\,
            sr => \N__20955\
        );

    \uu0.l_count_5_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__9037\,
            in1 => \_gnd_net_\,
            in2 => \N__9058\,
            in3 => \N__9097\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => \N__9073\,
            sr => \N__20955\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9053\,
            in2 => \_gnd_net_\,
            in3 => \N__9036\,
            lcout => \uu0.un88_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_2_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__13748\,
            in1 => \N__9378\,
            in2 => \N__9421\,
            in3 => \N__9405\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22292\,
            ce => \N__9767\,
            sr => \N__20957\
        );

    \buart.Z_rx.bitcount_es_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__9377\,
            in1 => \N__13749\,
            in2 => \N__10838\,
            in3 => \N__9461\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22292\,
            ce => \N__9767\,
            sr => \N__20957\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9568\,
            in2 => \_gnd_net_\,
            in3 => \N__9587\,
            lcout => \resetGen.un241_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9549\,
            lcout => \resetGen.reset_count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_RNILLLG7_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__9355\,
            in1 => \N__9348\,
            in2 => \_gnd_net_\,
            in3 => \N__9306\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15976\,
            in1 => \N__11149\,
            in2 => \_gnd_net_\,
            in3 => \N__21868\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__11833\,
            in1 => \N__9537\,
            in2 => \N__9574\,
            in3 => \N__9589\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__9534\,
            in1 => \N__9570\,
            in2 => \_gnd_net_\,
            in3 => \N__11832\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__11836\,
            in1 => \N__9510\,
            in2 => \N__9538\,
            in3 => \N__9232\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9588\,
            in1 => \N__9569\,
            in2 => \_gnd_net_\,
            in3 => \N__9495\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__11835\,
            in1 => \N__9536\,
            in2 => \N__9553\,
            in3 => \N__9550\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__11834\,
            in1 => \N__9535\,
            in2 => \N__9499\,
            in3 => \N__9511\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14797\,
            in2 => \_gnd_net_\,
            in3 => \N__21034\,
            lcout => \Lab_UT.didp.regrce2.LdAStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9735\,
            in1 => \N__9716\,
            in2 => \_gnd_net_\,
            in3 => \N__13752\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9672\,
            in1 => \N__9656\,
            in2 => \N__9606\,
            in3 => \N__9734\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9695\,
            in2 => \N__9481\,
            in3 => \N__9712\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9478\,
            in2 => \N__9469\,
            in3 => \N__9465\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__9682\,
            in1 => \N__9696\,
            in2 => \N__13764\,
            in3 => \N__9628\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__13751\,
            in1 => \_gnd_net_\,
            in2 => \N__9720\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__9657\,
            in1 => \N__9629\,
            in2 => \N__9643\,
            in3 => \N__13753\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__13750\,
            in1 => \N__13785\,
            in2 => \N__9631\,
            in3 => \N__18040\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9736\,
            in2 => \N__9721\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9697\,
            in2 => \_gnd_net_\,
            in3 => \N__9676\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13765\,
            in1 => \N__9673\,
            in2 => \_gnd_net_\,
            in3 => \N__9661\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__22273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9658\,
            in2 => \_gnd_net_\,
            in3 => \N__9634\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__9630\,
            in1 => \N__13758\,
            in2 => \N__9607\,
            in3 => \N__9610\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_3_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9927\,
            in1 => \N__9896\,
            in2 => \N__9831\,
            in3 => \N__10260\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__10228\,
            sr => \N__20948\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9845\,
            in2 => \_gnd_net_\,
            in3 => \N__9799\,
            lcout => OPEN,
            ltout => \uu2.vbuf_raddr.un448_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10165\,
            in1 => \N__9861\,
            in2 => \N__9868\,
            in3 => \N__9783\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__10228\,
            sr => \N__20948\
        );

    \uu2.r_addr_esr_7_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9784\,
            in1 => \N__9846\,
            in2 => \N__10171\,
            in3 => \N__9800\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__10228\,
            sr => \N__20948\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9926\,
            in1 => \N__9895\,
            in2 => \N__9830\,
            in3 => \N__10259\,
            lcout => \uu2.un404_ci_0\,
            ltout => \uu2.un404_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__10205\,
            in1 => \N__10117\,
            in2 => \N__9808\,
            in3 => \N__9801\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__10228\,
            sr => \N__20948\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10103\,
            in2 => \_gnd_net_\,
            in3 => \N__10204\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__13228\,
            in1 => \N__13108\,
            in2 => \N__11896\,
            in3 => \N__13177\,
            lcout => \uu2.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__21911\,
            in1 => \N__12810\,
            in2 => \N__10537\,
            in3 => \N__10741\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__9973\,
            in1 => \N__10699\,
            in2 => \_gnd_net_\,
            in3 => \N__21910\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__10512\,
            in1 => \N__10529\,
            in2 => \_gnd_net_\,
            in3 => \N__12808\,
            lcout => \uu2.N_34\,
            ltout => \uu2.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__10894\,
            in1 => \N__21913\,
            in2 => \N__9967\,
            in3 => \N__10566\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__10567\,
            in1 => \N__9946\,
            in2 => \N__21919\,
            in3 => \N__10783\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9945\,
            in1 => \N__10762\,
            in2 => \_gnd_net_\,
            in3 => \N__21909\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__10513\,
            in1 => \N__12809\,
            in2 => \N__10536\,
            in3 => \N__11148\,
            lcout => \uu2.N_31\,
            ltout => \uu2.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21912\,
            in2 => \N__9937\,
            in3 => \N__11713\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_2_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10140\,
            in1 => \N__9922\,
            in2 => \N__9900\,
            in3 => \N__10255\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => 'H',
            sr => \N__20941\
        );

    \uu2.r_addr_1_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10254\,
            in1 => \N__9891\,
            in2 => \_gnd_net_\,
            in3 => \N__10138\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => 'H',
            sr => \N__20941\
        );

    \uu2.r_addr_0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10253\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => 'H',
            sr => \N__20941\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10136\,
            in2 => \_gnd_net_\,
            in3 => \N__21036\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_4_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10197\,
            in1 => \N__10167\,
            in2 => \_gnd_net_\,
            in3 => \N__10139\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => 'H',
            sr => \N__20941\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11512\,
            in2 => \_gnd_net_\,
            in3 => \N__21885\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10642\,
            in2 => \_gnd_net_\,
            in3 => \N__10635\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_5_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10206\,
            in1 => \N__10166\,
            in2 => \N__10102\,
            in3 => \N__10141\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__20934\
        );

    \uu2.l_count_7_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10075\,
            in1 => \N__10001\,
            in2 => \N__10051\,
            in3 => \N__10033\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__20934\
        );

    \Lab_UT.didp.reset_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11206\,
            in1 => \_gnd_net_\,
            in2 => \N__12133\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__20934\
        );

    \Lab_UT.didp.ce_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12129\,
            in2 => \_gnd_net_\,
            in3 => \N__11205\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__20934\
        );

    \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14704\,
            in2 => \_gnd_net_\,
            in3 => \N__21033\,
            lcout => \Lab_UT.didp.regrce3.LdAMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10375\,
            in2 => \_gnd_net_\,
            in3 => \N__10339\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__17650\,
            in1 => \N__17688\,
            in2 => \_gnd_net_\,
            in3 => \N__14258\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17689\,
            in1 => \N__17312\,
            in2 => \N__10294\,
            in3 => \N__17763\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_3_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20521\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22302\,
            ce => \N__10291\,
            sr => \N__20932\
        );

    \Lab_UT.didp.regrce3.q_esr_0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14259\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22302\,
            ce => \N__10291\,
            sr => \N__20932\
        );

    \Lab_UT.didp.regrce3.q_esr_2_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20338\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22302\,
            ce => \N__10291\,
            sr => \N__20932\
        );

    \Lab_UT.didp.regrce3.q_esr_1_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20154\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22293\,
            ce => \N__10290\,
            sr => \N__20931\
        );

    \Lab_UT.alarmchar_latch_6_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011010"
        )
    port map (
            in0 => \N__11414\,
            in1 => \N__10270\,
            in2 => \N__11358\,
            in3 => \N__10501\,
            lcout => \G_184\,
            ltout => \G_184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__18364\,
            in1 => \_gnd_net_\,
            in2 => \N__10264\,
            in3 => \N__11575\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_idle_1_0_iclk_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__11348\,
            in1 => \N__11411\,
            in2 => \_gnd_net_\,
            in3 => \N__21035\,
            lcout => OPEN,
            ltout => \Lab_UT.un1_idle_1_0_iclkZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__10820\,
            in1 => \N__10915\,
            in2 => \N__10396\,
            in3 => \N__10479\,
            lcout => \G_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m59_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11410\,
            in1 => \N__12722\,
            in2 => \_gnd_net_\,
            in3 => \N__11347\,
            lcout => \Lab_UT.alarmstate_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11574\,
            in1 => \N__18363\,
            in2 => \_gnd_net_\,
            in3 => \N__10467\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__13638\,
            in1 => \N__11599\,
            in2 => \N__10393\,
            in3 => \N__11746\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11407\,
            in1 => \N__21023\,
            in2 => \_gnd_net_\,
            in3 => \N__11343\,
            lcout => \G_180\,
            ltout => \G_180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__11346\,
            in1 => \N__10500\,
            in2 => \N__10390\,
            in3 => \N__10951\,
            lcout => \G_181\,
            ltout => \G_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_0__m3_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__10942\,
            in1 => \N__12397\,
            in2 => \N__10387\,
            in3 => \N__11415\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__10384\,
            in1 => \N__11408\,
            in2 => \N__10378\,
            in3 => \N__10498\,
            lcout => \G_179\,
            ltout => \G_179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_armed_2_0_iso_i_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10504\,
            in3 => \N__11344\,
            lcout => \Lab_UT.un1_armed_2_0_iso_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_idle_5_0_iclk_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__11345\,
            in1 => \N__11409\,
            in2 => \_gnd_net_\,
            in3 => \N__10499\,
            lcout => OPEN,
            ltout => \Lab_UT.un1_idle_5_0_iclkZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__10468\,
            in1 => \N__10819\,
            in2 => \N__10483\,
            in3 => \N__10480\,
            lcout => \G_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20326\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22274\,
            ce => \N__15481\,
            sr => \N__20963\
        );

    \buart.Z_rx.shifter_0_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20110\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22271\,
            ce => \N__15480\,
            sr => \N__20965\
        );

    \buart.Z_tx.shifter_7_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21697\,
            in1 => \N__10423\,
            in2 => \_gnd_net_\,
            in3 => \N__10456\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => \N__21622\,
            sr => \N__20971\
        );

    \buart.Z_tx.shifter_8_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21696\,
            in2 => \_gnd_net_\,
            in3 => \N__10432\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => \N__21622\,
            sr => \N__20971\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15871\,
            in1 => \N__21867\,
            in2 => \_gnd_net_\,
            in3 => \N__13338\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__13516\,
            in1 => \N__13498\,
            in2 => \_gnd_net_\,
            in3 => \N__21021\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__21791\,
            in1 => \N__20682\,
            in2 => \_gnd_net_\,
            in3 => \N__13176\,
            lcout => \uu2.w_addr_displaying_RNI03P31Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__16153\,
            in1 => \N__11488\,
            in2 => \_gnd_net_\,
            in3 => \N__10795\,
            lcout => \uu2.un28_w_addr_user_i\,
            ltout => \uu2.un28_w_addr_user_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNID65PE_4_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10540\,
            in3 => \N__15822\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI43E87_4_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__16152\,
            in1 => \N__21020\,
            in2 => \_gnd_net_\,
            in3 => \N__10794\,
            lcout => \uu2.w_addr_user_RNI43E87Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIKIPH1_8_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20684\,
            in1 => \N__21782\,
            in2 => \N__16136\,
            in3 => \N__13342\,
            lcout => \uu2.un51_w_data_displaying_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11119\,
            in2 => \_gnd_net_\,
            in3 => \N__20683\,
            lcout => OPEN,
            ltout => \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIASLS1_8_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21781\,
            in1 => \N__16126\,
            in2 => \N__10516\,
            in3 => \N__13341\,
            lcout => \uu2.w_data_displaying_2_i_a2_i_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16127\,
            in1 => \N__20687\,
            in2 => \N__21792\,
            in3 => \N__11124\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__13253\,
            sr => \N__20895\
        );

    \uu2.w_addr_displaying_fast_nesr_3_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20685\,
            in1 => \N__21784\,
            in2 => \N__11135\,
            in3 => \N__11943\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__13253\,
            sr => \N__20895\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21783\,
            in1 => \N__20686\,
            in2 => \N__16468\,
            in3 => \N__11120\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__13253\,
            sr => \N__20895\
        );

    \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001000"
        )
    port map (
            in0 => \N__21780\,
            in1 => \N__12001\,
            in2 => \N__16135\,
            in3 => \N__11029\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0FGN6_4_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10585\,
            in2 => \N__10579\,
            in3 => \N__11059\,
            lcout => \uu2.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10648\,
            in1 => \N__10552\,
            in2 => \_gnd_net_\,
            in3 => \N__11014\,
            lcout => OPEN,
            ltout => \uu2.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__10576\,
            in1 => \N__10546\,
            in2 => \N__10570\,
            in3 => \N__12013\,
            lcout => \uu2.bitmap_pmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__16457\,
            in1 => \N__13339\,
            in2 => \_gnd_net_\,
            in3 => \N__12104\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNICM7R_180_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16780\,
            in1 => \N__12190\,
            in2 => \_gnd_net_\,
            in3 => \N__11947\,
            lcout => OPEN,
            ltout => \uu2.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__16458\,
            in1 => \N__16332\,
            in2 => \N__10558\,
            in3 => \N__12166\,
            lcout => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2\,
            ltout => \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__11049\,
            in1 => \N__10665\,
            in2 => \N__10555\,
            in3 => \N__16731\,
            lcout => \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__13340\,
            in1 => \N__11035\,
            in2 => \_gnd_net_\,
            in3 => \N__16333\,
            lcout => \uu2.bitmap_pmux_u_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__10666\,
            in1 => \N__16732\,
            in2 => \N__11053\,
            in3 => \N__10654\,
            lcout => \uu2.w_addr_displaying_RNI0NG56Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13809\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__20942\
        );

    \uu2.trig_rd_det_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10636\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__20942\
        );

    \uu2.trig_rd_det_0_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14357\,
            in2 => \_gnd_net_\,
            in3 => \N__14322\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__20942\
        );

    \buart.Z_rx.hh_0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10624\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__20942\
        );

    \uu0.sec_clkD_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13559\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0_sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22311\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11268\,
            in2 => \_gnd_net_\,
            in3 => \N__13558\,
            lcout => \oneSecStrb\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18260\,
            in1 => \N__18356\,
            in2 => \N__18455\,
            in3 => \N__12490\,
            lcout => \Lab_UT.dispString.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111110101111"
        )
    port map (
            in0 => \N__11487\,
            in1 => \N__11464\,
            in2 => \N__22357\,
            in3 => \N__11443\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14260\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22303\,
            ce => \N__12316\,
            sr => \N__20935\
        );

    \Lab_UT.didp.regrce4.q_esr_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20184\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22303\,
            ce => \N__12316\,
            sr => \N__20935\
        );

    \Lab_UT.didp.regrce4.q_esr_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20337\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22303\,
            ce => \N__12316\,
            sr => \N__20935\
        );

    \Lab_UT.didp.regrce4.q_esr_3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20522\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22303\,
            ce => \N__12316\,
            sr => \N__20935\
        );

    \Lab_UT.dispString.cnt_RNIH15E_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18426\,
            in1 => \N__18244\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dispString.un42_dOutP_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18350\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22294\,
            ce => 'H',
            sr => \N__20933\
        );

    \Lab_UT.dispString.cnt_0_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__18349\,
            in1 => \N__11657\,
            in2 => \N__18261\,
            in3 => \N__18427\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22294\,
            ce => 'H',
            sr => \N__20933\
        );

    \Lab_UT.didp.ce_0_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11656\,
            in1 => \N__17788\,
            in2 => \_gnd_net_\,
            in3 => \N__21287\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22294\,
            ce => 'H',
            sr => \N__20933\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__11774\,
            in1 => \N__12285\,
            in2 => \N__12604\,
            in3 => \N__14153\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11687\,
            in2 => \N__10669\,
            in3 => \N__17396\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10754\,
            in1 => \N__10886\,
            in2 => \_gnd_net_\,
            in3 => \N__11702\,
            lcout => \uu2.un1_w_user_crZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11703\,
            in1 => \N__10755\,
            in2 => \N__10698\,
            in3 => \N__10776\,
            lcout => OPEN,
            ltout => \uu2.un1_w_user_lfZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un20_w_addr_user_1_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__10717\,
            in1 => \N__11459\,
            in2 => \N__10798\,
            in3 => \N__11438\,
            lcout => \uu2.un20_w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_4_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__11504\,
            in1 => \N__10685\,
            in2 => \N__10740\,
            in3 => \N__10775\,
            lcout => \uu2.un1_w_user_crZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__18358\,
            in1 => \N__18267\,
            in2 => \_gnd_net_\,
            in3 => \N__10858\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_3_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__10887\,
            in1 => \_gnd_net_\,
            in2 => \N__11508\,
            in3 => \N__10733\,
            lcout => \uu2.un1_w_user_lfZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__18357\,
            in1 => \_gnd_net_\,
            in2 => \N__18448\,
            in3 => \N__18265\,
            lcout => \Lab_UT.dispString.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__18266\,
            in1 => \N__11776\,
            in2 => \N__10711\,
            in3 => \N__13361\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__11567\,
            in1 => \N__18362\,
            in2 => \N__11254\,
            in3 => \N__10870\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__18361\,
            in1 => \N__11566\,
            in2 => \N__11287\,
            in3 => \N__10914\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__10903\,
            in1 => \N__11747\,
            in2 => \N__10897\,
            in3 => \N__13424\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_0_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__11532\,
            in1 => \N__11353\,
            in2 => \N__21041\,
            in3 => \N__11413\,
            lcout => \G_186\,
            ltout => \G_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__18447\,
            in1 => \_gnd_net_\,
            in2 => \N__10873\,
            in3 => \N__18359\,
            lcout => \Lab_UT.dispString.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_4_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__10869\,
            in1 => \N__10977\,
            in2 => \N__21042\,
            in3 => \N__11354\,
            lcout => \G_187\,
            ltout => \G_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__11565\,
            in1 => \N__11250\,
            in2 => \N__10861\,
            in3 => \N__18360\,
            lcout => \Lab_UT.dispString.dOutP_1_iv_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001111"
        )
    port map (
            in0 => \N__10966\,
            in1 => \N__10941\,
            in2 => \N__10981\,
            in3 => \N__12396\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.justentered_latch_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__12395\,
            in1 => \N__10964\,
            in2 => \N__10852\,
            in3 => \N__21040\,
            lcout => \G_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11352\,
            in2 => \_gnd_net_\,
            in3 => \N__11412\,
            lcout => \G_182\,
            ltout => \G_182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__10965\,
            in1 => \N__10940\,
            in2 => \N__10954\,
            in3 => \N__12394\,
            lcout => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_7_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15378\,
            in1 => \N__15558\,
            in2 => \N__12956\,
            in3 => \N__12865\,
            lcout => \Lab_UT.dictrl.g1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_3_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15698\,
            in1 => \N__12933\,
            in2 => \N__20028\,
            in3 => \N__15377\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15553\,
            in1 => \N__12864\,
            in2 => \N__10945\,
            in3 => \N__19578\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__15699\,
            in1 => \_gnd_net_\,
            in2 => \N__20029\,
            in3 => \N__15554\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20127\,
            in1 => \N__11806\,
            in2 => \N__10927\,
            in3 => \N__15194\,
            lcout => \Lab_UT.dictrl.g1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__20441\,
            in1 => \N__20126\,
            in2 => \_gnd_net_\,
            in3 => \N__20303\,
            lcout => \Lab_UT.dictrl.g2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__12937\,
            in1 => \N__20442\,
            in2 => \N__15565\,
            in3 => \N__12866\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_5_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__11785\,
            in1 => \N__10924\,
            in2 => \N__10918\,
            in3 => \N__21439\,
            lcout => \Lab_UT.dictrl.N_55_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15563\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__15479\,
            sr => \N__20966\
        );

    \buart.Z_rx.shifter_4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12893\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__15479\,
            sr => \N__20966\
        );

    \buart.Z_rx.shifter_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12962\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__15479\,
            sr => \N__20966\
        );

    \buart.Z_rx.shifter_3_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15389\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__15479\,
            sr => \N__20966\
        );

    \buart.Z_rx.shifter_2_rep1_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20459\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22268\,
            ce => \N__15478\,
            sr => \N__20967\
        );

    \buart.Z_rx.shifter_3_rep2_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15390\,
            lcout => bu_rx_data_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22268\,
            ce => \N__15478\,
            sr => \N__20967\
        );

    \buart.Z_rx.shifter_fast_2_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20460\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22268\,
            ce => \N__15478\,
            sr => \N__20967\
        );

    \buart.Z_rx.shifter_fast_5_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12963\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22266\,
            ce => \N__15476\,
            sr => \N__20968\
        );

    \buart.Z_rx.shifter_0_rep1_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20155\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22266\,
            ce => \N__15476\,
            sr => \N__20968\
        );

    \buart.Z_rx.shifter_3_rep1_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15403\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22266\,
            ce => \N__15476\,
            sr => \N__20968\
        );

    \buart.Z_rx.shifter_fast_3_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15404\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => \N__15475\,
            sr => \N__20970\
        );

    \uu2.w_addr_user_2_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__21945\,
            in1 => \N__15966\,
            in2 => \N__20743\,
            in3 => \N__11000\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_user_1_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10998\,
            in1 => \N__15962\,
            in2 => \_gnd_net_\,
            in3 => \N__20738\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_user_0_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10997\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_user_4_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10999\,
            in1 => \N__15923\,
            in2 => \_gnd_net_\,
            in3 => \N__16185\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_user_5_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16186\,
            in1 => \N__15439\,
            in2 => \N__15928\,
            in3 => \N__11001\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_user_6_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11002\,
            in1 => \N__15927\,
            in2 => \N__15904\,
            in3 => \N__16051\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__15834\
        );

    \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21022\,
            in2 => \_gnd_net_\,
            in3 => \N__13932\,
            lcout => \uu2.N_33_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110111110"
        )
    port map (
            in0 => \N__13160\,
            in1 => \N__16251\,
            in2 => \N__16467\,
            in3 => \N__11987\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101000010"
        )
    port map (
            in0 => \N__11131\,
            in1 => \N__16119\,
            in2 => \N__11038\,
            in3 => \N__11028\,
            lcout => \uu2.bitmap_pmux_sn_i5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12097\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010010"
        )
    port map (
            in0 => \N__11988\,
            in1 => \N__16331\,
            in2 => \N__12106\,
            in3 => \N__16462\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16429\,
            in2 => \N__11017\,
            in3 => \N__11953\,
            lcout => \uu2.N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__12101\,
            in1 => \_gnd_net_\,
            in2 => \N__16262\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__13261\,
            sr => \N__20899\
        );

    \uu2.w_addr_displaying_fast_nesr_1_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16255\,
            in2 => \_gnd_net_\,
            in3 => \N__12102\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__13261\,
            sr => \N__20899\
        );

    \uu2.w_addr_displaying_nesr_1_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__12103\,
            in1 => \_gnd_net_\,
            in2 => \N__16263\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1_rep1_nesrC_net\,
            ce => \N__13261\,
            sr => \N__20899\
        );

    \uu2.bitmap_197_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__17374\,
            in1 => \N__16564\,
            in2 => \N__16387\,
            in3 => \N__16420\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20896\
        );

    \uu2.bitmap_RNITSCU1_69_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__11008\,
            in1 => \N__16345\,
            in2 => \N__11129\,
            in3 => \N__16513\,
            lcout => \uu2.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11110\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20896\
        );

    \uu2.w_addr_displaying_fast_2_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11112\,
            in1 => \N__13957\,
            in2 => \N__20703\,
            in3 => \N__11989\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20896\
        );

    \uu2.w_addr_displaying_2_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20681\,
            in1 => \N__11111\,
            in2 => \N__13960\,
            in3 => \N__21776\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__20896\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21775\,
            in1 => \N__16112\,
            in2 => \N__11130\,
            in3 => \N__20680\,
            lcout => \uu2.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000100000000"
        )
    port map (
            in0 => \N__16111\,
            in1 => \N__21774\,
            in2 => \N__11128\,
            in3 => \N__11848\,
            lcout => \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101000001000"
        )
    port map (
            in0 => \N__21773\,
            in1 => \N__20679\,
            in2 => \N__16128\,
            in3 => \N__13175\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12122\,
            in1 => \N__17142\,
            in2 => \_gnd_net_\,
            in3 => \N__11192\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => 'H',
            sr => \N__20945\
        );

    \Lab_UT.didp.ce_1_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13469\,
            in1 => \N__11169\,
            in2 => \N__11654\,
            in3 => \N__17604\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => 'H',
            sr => \N__20945\
        );

    \Lab_UT.didp.reset_0_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17605\,
            in1 => \N__13470\,
            in2 => \N__11173\,
            in3 => \N__11637\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => 'H',
            sr => \N__20945\
        );

    \Lab_UT.didp.reset_2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12123\,
            in1 => \N__17143\,
            in2 => \_gnd_net_\,
            in3 => \N__11193\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => 'H',
            sr => \N__20945\
        );

    \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13468\,
            in1 => \N__11168\,
            in2 => \N__11653\,
            in3 => \N__17603\,
            lcout => \Lab_UT.didp.ce_12_1\,
            ltout => \Lab_UT.didp.ce_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12121\,
            in1 => \_gnd_net_\,
            in2 => \N__11179\,
            in3 => \N__17141\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13849\,
            in1 => \N__17440\,
            in2 => \N__11176\,
            in3 => \N__17050\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => 'H',
            sr => \N__20945\
        );

    \Lab_UT.didp.ce_RNIBN0Q1_2_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11229\,
            in2 => \_gnd_net_\,
            in3 => \N__16956\,
            lcout => \Lab_UT.didp.un1_dicLdMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17717\,
            in2 => \_gnd_net_\,
            in3 => \N__17277\,
            lcout => \Lab_UT.didp.countrce1.ce_12_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17278\,
            in1 => \N__17721\,
            in2 => \_gnd_net_\,
            in3 => \N__17602\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__17646\,
            in1 => \N__13462\,
            in2 => \N__11158\,
            in3 => \N__20511\,
            lcout => \Lab_UT.didp.countrce1.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16994\,
            in2 => \_gnd_net_\,
            in3 => \N__17941\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__16955\,
            in1 => \N__20336\,
            in2 => \N__11155\,
            in3 => \N__17225\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17226\,
            in1 => \N__17992\,
            in2 => \N__11152\,
            in3 => \N__17952\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__16995\,
            in1 => \N__16954\,
            in2 => \_gnd_net_\,
            in3 => \N__14265\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__13463\,
            in1 => \N__17302\,
            in2 => \N__17764\,
            in3 => \N__11296\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__13425\,
            in1 => \N__17045\,
            in2 => \N__13464\,
            in3 => \N__13826\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_3_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__13827\,
            in1 => \N__11686\,
            in2 => \N__11655\,
            in3 => \N__18433\,
            lcout => \Lab_UT.dispString.N_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18248\,
            in2 => \_gnd_net_\,
            in3 => \N__18319\,
            lcout => \Lab_UT.dispString.N_143\,
            ltout => \Lab_UT.dispString.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIKUO21_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__13564\,
            in2 => \N__11257\,
            in3 => \N__18432\,
            lcout => \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18434\,
            in1 => \N__11641\,
            in2 => \N__18268\,
            in3 => \N__18320\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000001"
        )
    port map (
            in0 => \N__16957\,
            in1 => \N__11233\,
            in2 => \N__18013\,
            in3 => \N__11212\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__16996\,
            in1 => \N__14438\,
            in2 => \N__12226\,
            in3 => \N__13871\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18242\,
            lcout => \Lab_UT.dispString.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIKUO21_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000101"
        )
    port map (
            in0 => \N__18243\,
            in1 => \N__18417\,
            in2 => \N__11665\,
            in3 => \N__18325\,
            lcout => \Lab_UT.dispString.N_102\,
            ltout => \Lab_UT.dispString.N_102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__18326\,
            in1 => \N__11573\,
            in2 => \N__11539\,
            in3 => \N__11536\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__11748\,
            in1 => \N__11521\,
            in2 => \N__11515\,
            in3 => \N__14400\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__11477\,
            in1 => \N__11460\,
            in2 => \_gnd_net_\,
            in3 => \N__11439\,
            lcout => \uu2.un4_w_user_data_rdyZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIFV4E_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18416\,
            in2 => \_gnd_net_\,
            in3 => \N__18324\,
            lcout => \Lab_UT.dispString.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNIHGGI1_3_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__17121\,
            in1 => \_gnd_net_\,
            in2 => \N__12339\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.un1_dicLdMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000010"
        )
    port map (
            in0 => \N__11422\,
            in1 => \N__17188\,
            in2 => \N__11365\,
            in3 => \N__13372\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__17728\,
            in1 => \N__11305\,
            in2 => \N__11299\,
            in3 => \N__13392\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__11775\,
            in1 => \N__12225\,
            in2 => \N__13879\,
            in3 => \N__11688\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__12603\,
            in1 => \N__11758\,
            in2 => \N__11752\,
            in3 => \N__12368\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__11749\,
            in1 => \N__11722\,
            in2 => \N__11716\,
            in3 => \N__13391\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__11689\,
            in1 => \N__12580\,
            in2 => \N__11664\,
            in3 => \N__16590\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14253\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22272\,
            ce => \N__11587\,
            sr => \N__20936\
        );

    \Lab_UT.didp.regrce2.q_esr_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20169\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22272\,
            ce => \N__11587\,
            sr => \N__20936\
        );

    \Lab_UT.didp.regrce2.q_esr_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20325\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22272\,
            ce => \N__11587\,
            sr => \N__20936\
        );

    \Lab_UT.didp.regrce2.q_esr_3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20487\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22272\,
            ce => \N__11587\,
            sr => \N__20936\
        );

    \Lab_UT.didp.regrce1.q_esr_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14257\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22270\,
            ce => \N__12574\,
            sr => \N__20938\
        );

    \Lab_UT.dictrl.g1_8_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19457\,
            in1 => \N__19735\,
            in2 => \N__15785\,
            in3 => \N__15708\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21438\,
            in1 => \N__11800\,
            in2 => \N__11791\,
            in3 => \N__19905\,
            lcout => \Lab_UT.dictrl.G_14_0_a2_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__19906\,
            in1 => \N__21437\,
            in2 => \_gnd_net_\,
            in3 => \N__12952\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_25_i_o3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__20312\,
            in1 => \N__20452\,
            in2 => \N__11788\,
            in3 => \N__20177\,
            lcout => \Lab_UT.dictrl.G_25_i_o3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__20311\,
            in1 => \N__20631\,
            in2 => \N__20162\,
            in3 => \N__15388\,
            lcout => \Lab_UT.dictrl.g0_5_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_6_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12883\,
            in2 => \_gnd_net_\,
            in3 => \N__12951\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20632\,
            in1 => \N__15564\,
            in2 => \N__11779\,
            in3 => \N__15387\,
            lcout => \Lab_UT.dictrl.g0_6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m37_N_2L1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14219\,
            in1 => \N__12867\,
            in2 => \N__20301\,
            in3 => \N__19991\,
            lcout => \Lab_UT.dictrl.m37_N_2LZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20261\,
            in2 => \_gnd_net_\,
            in3 => \N__14220\,
            lcout => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12990\,
            in2 => \_gnd_net_\,
            in3 => \N__13022\,
            lcout => \Lab_UT.dictrl.m13_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_4_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15386\,
            in1 => \N__20183\,
            in2 => \N__20483\,
            in3 => \N__14221\,
            lcout => OPEN,
            ltout => \resetGen.escKeyZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11812\,
            in2 => \N__11839\,
            in3 => \N__18078\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15561\,
            in1 => \N__12950\,
            in2 => \N__12885\,
            in3 => \N__20262\,
            lcout => \resetGen.escKeyZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_5_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__12949\,
            in1 => \N__12868\,
            in2 => \N__15787\,
            in3 => \N__15384\,
            lcout => \Lab_UT.dictrl.g1_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_5_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__15385\,
            in1 => \N__15562\,
            in2 => \N__21289\,
            in3 => \N__12884\,
            lcout => \Lab_UT.dictrl.G_25_i_o3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__19990\,
            in1 => \N__13028\,
            in2 => \N__19920\,
            in3 => \N__12992\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20274\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22265\,
            ce => \N__15477\,
            sr => \N__20969\
        );

    \buart.Z_rx.shifter_1_rep1_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22265\,
            ce => \N__15477\,
            sr => \N__20969\
        );

    \buart.Z_rx.shifter_2_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20461\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22265\,
            ce => \N__15477\,
            sr => \N__20969\
        );

    \Lab_UT.dictrl.g1_1_5_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13024\,
            in1 => \N__11910\,
            in2 => \N__15327\,
            in3 => \N__15646\,
            lcout => \Lab_UT.dictrl.g1_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12825\,
            in1 => \N__14689\,
            in2 => \N__11911\,
            in3 => \N__13023\,
            lcout => \Lab_UT.dictrl.g1_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m34_1_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12991\,
            in2 => \_gnd_net_\,
            in3 => \N__15645\,
            lcout => \Lab_UT.dictrl.m34Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_8_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000100"
        )
    port map (
            in0 => \N__12796\,
            in1 => \N__13947\,
            in2 => \N__11895\,
            in3 => \N__16759\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20902\
        );

    \uu2.w_addr_displaying_8_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__13945\,
            in1 => \N__13312\,
            in2 => \N__12811\,
            in3 => \N__11886\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20902\
        );

    \uu2.w_addr_displaying_RNI0ES07_8_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011111111"
        )
    port map (
            in0 => \N__13311\,
            in1 => \N__12804\,
            in2 => \N__11893\,
            in3 => \N__21866\,
            lcout => \uu2.w_addr_displaying_RNI0ES07Z0Z_8\,
            ltout => \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11882\,
            in2 => \N__11899\,
            in3 => \N__13173\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20902\
        );

    \uu2.w_addr_displaying_5_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__13174\,
            in1 => \N__13946\,
            in2 => \N__11894\,
            in3 => \N__13102\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_8C_net\,
            ce => 'H',
            sr => \N__20902\
        );

    \uu2.w_addr_displaying_ness_RNO_0_6_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__13101\,
            in1 => \N__11881\,
            in2 => \_gnd_net_\,
            in3 => \N__13172\,
            lcout => \uu2.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000011000"
        )
    port map (
            in0 => \N__13214\,
            in1 => \N__16311\,
            in2 => \N__13326\,
            in3 => \N__13099\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__13100\,
            in1 => \N__13310\,
            in2 => \N__16325\,
            in3 => \N__13215\,
            lcout => \uu2.bitmap_pmux_sn_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__14667\,
            in1 => \N__14502\,
            in2 => \N__14628\,
            in3 => \N__14576\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__20901\
        );

    \uu2.bitmap_75_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__14577\,
            in1 => \N__14621\,
            in2 => \N__14506\,
            in3 => \N__14668\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__20901\
        );

    \uu2.bitmap_203_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__14666\,
            in1 => \N__14501\,
            in2 => \N__14627\,
            in3 => \N__14575\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__20901\
        );

    \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__11986\,
            in1 => \N__11945\,
            in2 => \_gnd_net_\,
            in3 => \N__11968\,
            lcout => \uu2.bitmap_pmux_sn_N_54_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIJS4P_162_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11946\,
            in1 => \N__16501\,
            in2 => \_gnd_net_\,
            in3 => \N__13477\,
            lcout => OPEN,
            ltout => \uu2.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13522\,
            in2 => \N__11962\,
            in3 => \N__11959\,
            lcout => \uu2.bitmap_RNI2Q8F1Z0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIBPBO_40_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__11944\,
            in1 => \N__11917\,
            in2 => \N__13486\,
            in3 => \N__16761\,
            lcout => \uu2.bitmap_pmux_26_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011100011111"
        )
    port map (
            in0 => \N__16835\,
            in1 => \N__16881\,
            in2 => \N__16810\,
            in3 => \N__16912\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__20900\
        );

    \uu2.bitmap_221_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__16911\,
            in1 => \N__16806\,
            in2 => \N__16885\,
            in3 => \N__16834\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__20900\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12105\,
            lcout => \uu2.N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI6MCU1_93_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__16236\,
            in2 => \N__12067\,
            in3 => \N__16198\,
            lcout => \uu2.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIPIHG1_75_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__16235\,
            in1 => \N__12055\,
            in2 => \N__12049\,
            in3 => \N__13969\,
            lcout => OPEN,
            ltout => \uu2.N_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__16138\,
            in1 => \N__12036\,
            in2 => \N__12040\,
            in3 => \N__12139\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_27_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI72CH8_69_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__12037\,
            in1 => \N__12028\,
            in2 => \N__12022\,
            in3 => \N__12019\,
            lcout => \uu2.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__14025\,
            in1 => \N__14062\,
            in2 => \N__14131\,
            in3 => \N__14091\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_212_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__14090\,
            in1 => \N__14117\,
            in2 => \N__14068\,
            in3 => \N__14024\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_84_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__14027\,
            in1 => \N__14064\,
            in2 => \N__14133\,
            in3 => \N__14093\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_180_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__14089\,
            in1 => \N__14116\,
            in2 => \N__14067\,
            in3 => \N__14023\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_52_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__14026\,
            in1 => \N__14063\,
            in2 => \N__14132\,
            in3 => \N__14092\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_RNIB3QK_52_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__12178\,
            in2 => \_gnd_net_\,
            in3 => \N__12172\,
            lcout => \uu2.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__14028\,
            in1 => \N__14065\,
            in2 => \N__14134\,
            in3 => \N__14094\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__20897\
        );

    \uu2.bitmap_RNIRMQA1_84_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__12154\,
            in1 => \N__13990\,
            in2 => \N__12148\,
            in3 => \N__16717\,
            lcout => \uu2.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13602\,
            in1 => \N__14297\,
            in2 => \N__12256\,
            in3 => \N__12457\,
            lcout => \Lab_UT.didp.un24_ce_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001101"
        )
    port map (
            in0 => \N__17889\,
            in1 => \N__16671\,
            in2 => \N__12523\,
            in3 => \N__14164\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__14296\,
            in2 => \_gnd_net_\,
            in3 => \N__12373\,
            lcout => \Lab_UT.sec1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__13570\,
            in1 => \N__20339\,
            in2 => \N__17895\,
            in3 => \N__12253\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__12254\,
            in1 => \N__12519\,
            in2 => \N__12301\,
            in3 => \N__16650\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12286\,
            in1 => \N__12248\,
            in2 => \_gnd_net_\,
            in3 => \N__17521\,
            lcout => \Lab_UT.sec1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17519\,
            in1 => \N__12456\,
            in2 => \_gnd_net_\,
            in3 => \N__12489\,
            lcout => \Lab_UT.sec1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__14298\,
            in1 => \N__12252\,
            in2 => \_gnd_net_\,
            in3 => \N__13601\,
            lcout => \Lab_UT.didp.countrce2.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__12298\,
            in1 => \N__20523\,
            in2 => \N__17896\,
            in3 => \N__12458\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__16657\,
            in1 => \N__12459\,
            in2 => \N__12289\,
            in3 => \N__12517\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17578\,
            in1 => \N__12281\,
            in2 => \N__12255\,
            in3 => \N__13631\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17397\,
            in1 => \N__14532\,
            in2 => \N__17940\,
            in3 => \N__17429\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__12224\,
            in2 => \_gnd_net_\,
            in3 => \N__17510\,
            lcout => \Lab_UT.min2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101010101"
        )
    port map (
            in0 => \N__20187\,
            in1 => \N__14301\,
            in2 => \N__13609\,
            in3 => \N__17894\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__12518\,
            in1 => \N__13606\,
            in2 => \N__12493\,
            in3 => \N__16656\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13662\,
            in1 => \N__12482\,
            in2 => \N__12460\,
            in3 => \N__13595\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14374\,
            in1 => \N__12430\,
            in2 => \N__12424\,
            in3 => \N__12421\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12349\,
            in1 => \N__12415\,
            in2 => \N__12406\,
            in3 => \N__12403\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__12369\,
            in1 => \N__17227\,
            in2 => \N__14305\,
            in3 => \N__14154\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__17109\,
            in1 => \N__14437\,
            in2 => \_gnd_net_\,
            in3 => \N__14264\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000001"
        )
    port map (
            in0 => \N__14746\,
            in1 => \N__17110\,
            in2 => \N__12343\,
            in3 => \N__12340\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__21251\,
            in1 => \N__20615\,
            in2 => \N__18949\,
            in3 => \N__21025\,
            lcout => \Lab_UT.didp.regrce4.LdAMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18368\,
            in1 => \N__18252\,
            in2 => \N__18456\,
            in3 => \N__14531\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__18369\,
            in2 => \N__12583\,
            in3 => \N__13661\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14809\,
            in2 => \_gnd_net_\,
            in3 => \N__21024\,
            lcout => \Lab_UT.didp.regrce1.LdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20170\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__12567\,
            sr => \N__20939\
        );

    \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20330\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__12567\,
            sr => \N__20939\
        );

    \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20515\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__12567\,
            sr => \N__20939\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__19053\,
            in1 => \N__15223\,
            in2 => \N__15198\,
            in3 => \N__13048\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000001111"
        )
    port map (
            in0 => \N__12547\,
            in1 => \N__12535\,
            in2 => \N__12529\,
            in3 => \N__21166\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__19258\,
            in1 => \N__18066\,
            in2 => \N__12526\,
            in3 => \N__12637\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_25_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__18157\,
            in1 => \N__17824\,
            in2 => \N__12640\,
            in3 => \N__12631\,
            lcout => \Lab_UT.un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__19256\,
            in1 => \N__18065\,
            in2 => \N__18741\,
            in3 => \N__12724\,
            lcout => \Lab_UT.dictrl.G_25_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__21167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19052\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__18067\,
            in1 => \N__19257\,
            in2 => \N__18601\,
            in3 => \N__21058\,
            lcout => \Lab_UT.dictrl.G_25_i_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__19822\,
            in1 => \N__20037\,
            in2 => \N__19919\,
            in3 => \N__19588\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_18_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__12646\,
            in2 => \N__12625\,
            in3 => \N__21429\,
            lcout => \Lab_UT.dictrl.N_22_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__21428\,
            in1 => \N__15186\,
            in2 => \N__18770\,
            in3 => \N__19636\,
            lcout => \Lab_UT.dictrl.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__12673\,
            in1 => \N__12622\,
            in2 => \N__12616\,
            in3 => \N__21430\,
            lcout => \Lab_UT.dictrl.N_57_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__19455\,
            in1 => \N__19731\,
            in2 => \_gnd_net_\,
            in3 => \N__15788\,
            lcout => \shifter_1_rep1_RNI0FPF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__15789\,
            in1 => \N__19821\,
            in2 => \N__19738\,
            in3 => \N__19456\,
            lcout => \N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001100110"
        )
    port map (
            in0 => \N__21427\,
            in1 => \N__12661\,
            in2 => \N__18769\,
            in3 => \N__21159\,
            lcout => \Lab_UT.dictrl.m19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18046\,
            in1 => \N__12772\,
            in2 => \N__19245\,
            in3 => \N__12715\,
            lcout => \Lab_UT.didp.g0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19908\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15259\,
            in1 => \N__20469\,
            in2 => \N__12676\,
            in3 => \N__12740\,
            lcout => \Lab_UT.dictrl.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12667\,
            lcout => \Lab_UT.dictrl.N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__19907\,
            in1 => \N__13039\,
            in2 => \N__19723\,
            in3 => \N__12994\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__19820\,
            in1 => \_gnd_net_\,
            in2 => \N__12655\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m37_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__12652\,
            in2 => \N__15307\,
            in3 => \N__12957\,
            lcout => \Lab_UT.dictrl.next_state6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_8_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14222\,
            in1 => \N__15258\,
            in2 => \N__12742\,
            in3 => \N__20033\,
            lcout => \Lab_UT.dictrl.N_72_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m34_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15560\,
            in1 => \N__12886\,
            in2 => \N__15306\,
            in3 => \N__12958\,
            lcout => \Lab_UT.dictrl.N_67_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110101010"
        )
    port map (
            in0 => \N__12748\,
            in1 => \N__12741\,
            in2 => \N__15257\,
            in3 => \N__12763\,
            lcout => OPEN,
            ltout => \Lab_UT.i8_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_2_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12754\,
            in2 => \N__12775\,
            in3 => \N__21168\,
            lcout => \Lab_UT.didp.g0_0_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15225\,
            in1 => \N__20014\,
            in2 => \N__15715\,
            in3 => \N__15184\,
            lcout => \Lab_UT.dictrl.g0_0_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__21278\,
            in2 => \_gnd_net_\,
            in3 => \N__21419\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__19800\,
            in1 => \N__20015\,
            in2 => \N__12757\,
            in3 => \N__19587\,
            lcout => \Lab_UT.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__19070\,
            in2 => \_gnd_net_\,
            in3 => \N__15224\,
            lcout => \Lab_UT.dictrl.g0_0_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21169\,
            in1 => \N__15185\,
            in2 => \N__21440\,
            in3 => \N__21288\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15783\,
            in2 => \_gnd_net_\,
            in3 => \N__19451\,
            lcout => \Lab_UT.dictrl.m22Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__19695\,
            in1 => \N__15786\,
            in2 => \_gnd_net_\,
            in3 => \N__19452\,
            lcout => \Lab_UT.dictrl.gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m5_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__12826\,
            in1 => \N__19365\,
            in2 => \N__19494\,
            in3 => \N__15649\,
            lcout => \N_63_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15624\,
            in2 => \_gnd_net_\,
            in3 => \N__19403\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_10_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15076\,
            in1 => \N__19453\,
            in2 => \N__13051\,
            in3 => \N__12894\,
            lcout => \Lab_UT.dictrl.N_72_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m7_a0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13038\,
            in2 => \_gnd_net_\,
            in3 => \N__12993\,
            lcout => m7_a0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_rep1_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12964\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__15473\,
            sr => \N__20972\
        );

    \buart.Z_rx.shifter_fast_4_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_fast_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__15473\,
            sr => \N__20972\
        );

    \buart.Z_rx.shifter_fast_6_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__15473\,
            sr => \N__20972\
        );

    \buart.Z_rx.shifter_fast_7_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15599\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22264\,
            ce => \N__15473\,
            sr => \N__20972\
        );

    \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__16321\,
            in1 => \N__13103\,
            in2 => \N__13224\,
            in3 => \N__13170\,
            lcout => \uu2.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_6_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100000001111"
        )
    port map (
            in0 => \N__13325\,
            in1 => \N__16323\,
            in2 => \N__13270\,
            in3 => \N__13220\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_ness_6C_net\,
            ce => \N__13260\,
            sr => \N__20905\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13219\,
            in1 => \N__16047\,
            in2 => \_gnd_net_\,
            in3 => \N__21901\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13171\,
            in1 => \N__16187\,
            in2 => \_gnd_net_\,
            in3 => \N__21899\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21900\,
            in1 => \N__15443\,
            in2 => \_gnd_net_\,
            in3 => \N__13104\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__15444\,
            in1 => \N__16188\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.un426_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16322\,
            in1 => \N__16013\,
            in2 => \_gnd_net_\,
            in3 => \N__21902\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16050\,
            lcout => \uu2.vbuf_w_addr_user.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13943\,
            in1 => \N__13896\,
            in2 => \_gnd_net_\,
            in3 => \N__16324\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.w_addr_displaying_0_rep1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13944\,
            in2 => \_gnd_net_\,
            in3 => \N__16249\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.bitmap_111_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13563\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.vram_rd_clk_det_0_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14362\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.vram_rd_clk_det_1_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13512\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.bitmap_296_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__14584\,
            in1 => \N__14609\,
            in2 => \N__14500\,
            in3 => \N__14658\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \uu2.bitmap_168_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__14657\,
            in1 => \N__14488\,
            in2 => \N__14622\,
            in3 => \N__14583\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7C_net\,
            ce => 'H',
            sr => \N__20903\
        );

    \Lab_UT.dictrl.next_state_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011000000"
        )
    port map (
            in0 => \N__18661\,
            in1 => \N__21282\,
            in2 => \N__18634\,
            in3 => \N__21165\,
            lcout => \Lab_UT.dictrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22333\,
            ce => \N__19342\,
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__13471\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \Lab_UT.sec2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17725\,
            in1 => \N__13393\,
            in2 => \_gnd_net_\,
            in3 => \N__17508\,
            lcout => \Lab_UT.sec2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17505\,
            in1 => \_gnd_net_\,
            in2 => \N__17180\,
            in3 => \N__13371\,
            lcout => \Lab_UT.min2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14451\,
            in1 => \N__13878\,
            in2 => \_gnd_net_\,
            in3 => \N__17507\,
            lcout => \Lab_UT.min1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14452\,
            in2 => \_gnd_net_\,
            in3 => \N__16636\,
            lcout => \Lab_UT.didp.reset_12_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13837\,
            in1 => \N__17046\,
            in2 => \_gnd_net_\,
            in3 => \N__17506\,
            lcout => \Lab_UT.min1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13813\,
            in1 => \N__15585\,
            in2 => \_gnd_net_\,
            in3 => \N__13795\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13669\,
            in1 => \N__13607\,
            in2 => \_gnd_net_\,
            in3 => \N__17503\,
            lcout => \Lab_UT.sec1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17502\,
            in1 => \N__17591\,
            in2 => \_gnd_net_\,
            in3 => \N__13639\,
            lcout => \Lab_UT.sec2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16635\,
            in2 => \_gnd_net_\,
            in3 => \N__14450\,
            lcout => \Lab_UT.didp.countrce4.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__13608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14299\,
            lcout => \Lab_UT.didp.countrce2.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14401\,
            in1 => \N__17271\,
            in2 => \_gnd_net_\,
            in3 => \N__17504\,
            lcout => \Lab_UT.sec2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__14358\,
            in1 => \N__14326\,
            in2 => \N__21043\,
            in3 => \N__21657\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__14300\,
            in1 => \N__17890\,
            in2 => \_gnd_net_\,
            in3 => \N__14266\,
            lcout => \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17501\,
            in1 => \N__17235\,
            in2 => \_gnd_net_\,
            in3 => \N__14158\,
            lcout => \Lab_UT.min2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__14130\,
            in1 => \N__14095\,
            in2 => \N__14066\,
            in3 => \N__14029\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20898\
        );

    \uu2.bitmap_RNIOPSS_212_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__14002\,
            in1 => \N__13996\,
            in2 => \N__13984\,
            in3 => \N__16714\,
            lcout => \uu2.bitmap_pmux_17_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13958\,
            in2 => \_gnd_net_\,
            in3 => \N__13983\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20898\
        );

    \uu2.bitmap_RNI65TM_72_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__13982\,
            in1 => \N__14674\,
            in2 => \N__14545\,
            in3 => \N__16715\,
            lcout => \uu2.bitmap_pmux_16_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_7_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__16716\,
            in1 => \N__13959\,
            in2 => \_gnd_net_\,
            in3 => \N__13900\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20898\
        );

    \uu2.bitmap_72_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__14564\,
            in1 => \N__14626\,
            in2 => \N__14499\,
            in3 => \N__14648\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20898\
        );

    \uu2.bitmap_200_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__14647\,
            in1 => \N__14484\,
            in2 => \N__14629\,
            in3 => \N__14563\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__20898\
        );

    \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17929\,
            in1 => \N__17500\,
            in2 => \_gnd_net_\,
            in3 => \N__14536\,
            lcout => \Lab_UT.min2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__16632\,
            in1 => \N__14433\,
            in2 => \N__17125\,
            in3 => \N__20199\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__14747\,
            in1 => \N__14773\,
            in2 => \N__14455\,
            in3 => \N__16633\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16631\,
            in1 => \N__14432\,
            in2 => \_gnd_net_\,
            in3 => \N__17431\,
            lcout => \Lab_UT.didp.countrce4.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__17044\,
            in1 => \N__17008\,
            in2 => \N__14754\,
            in3 => \N__14772\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__17762\,
            in1 => \N__17542\,
            in2 => \N__17319\,
            in3 => \N__17590\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__14396\,
            in1 => \N__16586\,
            in2 => \N__16634\,
            in3 => \N__17262\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__14771\,
            in1 => \N__16519\,
            in2 => \N__14755\,
            in3 => \N__17432\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20624\,
            in1 => \N__21376\,
            in2 => \N__21277\,
            in3 => \N__21135\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18079\,
            in2 => \_gnd_net_\,
            in3 => \N__21032\,
            lcout => \Lab_UT.bu_rx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__18119\,
            in1 => \N__17825\,
            in2 => \N__18087\,
            in3 => \N__14713\,
            lcout => \Lab_UT.dictrl.dicLdAMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22305\,
            ce => 'H',
            sr => \N__20943\
        );

    \Lab_UT.dictrl.state_ret_5_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__17826\,
            in1 => \N__18159\,
            in2 => \N__14824\,
            in3 => \N__18083\,
            lcout => \Lab_UT.dictrl.dicRun_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22305\,
            ce => 'H',
            sr => \N__20943\
        );

    \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21255\,
            in1 => \N__21375\,
            in2 => \_gnd_net_\,
            in3 => \N__14712\,
            lcout => \Lab_UT.LdAMones\,
            ltout => \Lab_UT.LdAMones_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14790\,
            in1 => \N__14808\,
            in2 => \N__14692\,
            in3 => \N__18463\,
            lcout => \Lab_UT.loadalarm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001010111"
        )
    port map (
            in0 => \N__19137\,
            in1 => \N__19267\,
            in2 => \N__18700\,
            in3 => \N__15087\,
            lcout => \Lab_UT.dictrl.state_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__18530\,
            sr => \N__20937\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000111111101"
        )
    port map (
            in0 => \N__15088\,
            in1 => \N__18699\,
            in2 => \N__19275\,
            in3 => \N__19138\,
            lcout => \Lab_UT.dictrl.state_ret_2_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__18530\,
            sr => \N__20937\
        );

    \Lab_UT.dictrl.state_ret_6_ess_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000111111101"
        )
    port map (
            in0 => \N__14872\,
            in1 => \N__19054\,
            in2 => \N__19276\,
            in3 => \N__14848\,
            lcout => \Lab_UT.dictrl.state_i_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__18530\,
            sr => \N__20937\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18486\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \Lab_UT.dictrl.m19_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_esr_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19266\,
            in1 => \N__18886\,
            in2 => \N__18745\,
            in3 => \N__18158\,
            lcout => \Lab_UT.dictrl.next_state66_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__18530\,
            sr => \N__20937\
        );

    \Lab_UT.dictrl.state_ret_5_RNICG571_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14820\,
            in1 => \N__21226\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \Lab_UT.LdASones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15007\,
            in1 => \N__15046\,
            in2 => \N__14973\,
            in3 => \N__18814\,
            lcout => \Lab_UT.next_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18817\,
            in1 => \N__14972\,
            in2 => \N__15055\,
            in3 => \N__15010\,
            lcout => \Lab_UT.dictrl.state_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15008\,
            in1 => \N__15047\,
            in2 => \N__14974\,
            in3 => \N__18815\,
            lcout => \Lab_UT.dictrl.state_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18816\,
            in1 => \N__14971\,
            in2 => \N__15054\,
            in3 => \N__15009\,
            lcout => \Lab_UT.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21225\,
            in1 => \N__20582\,
            in2 => \N__18559\,
            in3 => \N__21359\,
            lcout => \Lab_UT.LdAStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__18879\,
            in1 => \N__18733\,
            in2 => \_gnd_net_\,
            in3 => \N__19227\,
            lcout => \Lab_UT.state_i_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19226\,
            in2 => \N__18740\,
            in3 => \N__18878\,
            lcout => \Lab_UT.dictrl.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__14867\,
            in1 => \N__14844\,
            in2 => \N__19071\,
            in3 => \N__19228\,
            lcout => \Lab_UT_dictrl_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => \N__18538\,
            sr => \N__20944\
        );

    \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__19246\,
            in1 => \N__14943\,
            in2 => \N__14932\,
            in3 => \N__18560\,
            lcout => \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__18562\,
            in1 => \N__19051\,
            in2 => \N__14871\,
            in3 => \N__14944\,
            lcout => \Lab_UT.dictrl.next_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22281\,
            ce => \N__19331\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__14904\,
            in1 => \N__14892\,
            in2 => \N__15031\,
            in3 => \N__20613\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_20_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__18561\,
            in1 => \N__19049\,
            in2 => \N__14923\,
            in3 => \N__14920\,
            lcout => OPEN,
            ltout => \Lab_UT.next_state_1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.g0_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__18124\,
            in1 => \N__14914\,
            in2 => \N__14908\,
            in3 => \N__17809\,
            lcout => \Lab_UT.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__14905\,
            in1 => \N__14893\,
            in2 => \N__14884\,
            in3 => \N__20614\,
            lcout => \Lab_UT.dictrl.N_20\,
            ltout => \Lab_UT.dictrl.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__19244\,
            in1 => \N__14843\,
            in2 => \N__14827\,
            in3 => \N__19050\,
            lcout => \Lab_UT.next_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__20310\,
            in1 => \N__19827\,
            in2 => \N__20185\,
            in3 => \N__20030\,
            lcout => \N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__18840\,
            in2 => \N__19294\,
            in3 => \N__15064\,
            lcout => \Lab_UT.dictrl.G_14_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18487\,
            in2 => \_gnd_net_\,
            in3 => \N__21143\,
            lcout => \Lab_UT.dictrl.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__19828\,
            in1 => \N__19894\,
            in2 => \N__15022\,
            in3 => \N__21425\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__18841\,
            in1 => \N__20621\,
            in2 => \N__15013\,
            in3 => \N__14982\,
            lcout => \Lab_UT.dictrl.G_14_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19208\,
            in1 => \N__19061\,
            in2 => \_gnd_net_\,
            in3 => \N__18936\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_14_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011010000"
        )
    port map (
            in0 => \N__20616\,
            in1 => \N__14992\,
            in2 => \N__14986\,
            in3 => \N__14983\,
            lcout => \Lab_UT.dictrl.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111101"
        )
    port map (
            in0 => \N__19816\,
            in1 => \N__19121\,
            in2 => \N__19730\,
            in3 => \N__19869\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19713\,
            in1 => \N__15070\,
            in2 => \N__14947\,
            in3 => \N__19590\,
            lcout => \Lab_UT.dictrl.N_60_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__19062\,
            in1 => \N__15226\,
            in2 => \N__15199\,
            in3 => \N__19631\,
            lcout => \Lab_UT.dictrl.i8_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__19122\,
            in1 => \N__20468\,
            in2 => \_gnd_net_\,
            in3 => \N__19817\,
            lcout => OPEN,
            ltout => \N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001000"
        )
    port map (
            in0 => \N__19063\,
            in1 => \N__18948\,
            in2 => \N__15133\,
            in3 => \N__20622\,
            lcout => \Lab_UT.dictrl.G_6_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_5_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110100111"
        )
    port map (
            in0 => \N__21423\,
            in1 => \N__19818\,
            in2 => \N__20038\,
            in3 => \N__19589\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_3_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111111"
        )
    port map (
            in0 => \N__15130\,
            in1 => \N__15114\,
            in2 => \N__15118\,
            in3 => \N__21424\,
            lcout => \Lab_UT.dictrl.i9_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20623\,
            in1 => \N__19064\,
            in2 => \N__15661\,
            in3 => \N__15115\,
            lcout => \Lab_UT.dictrl.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__15103\,
            in1 => \N__15094\,
            in2 => \_gnd_net_\,
            in3 => \N__19090\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15711\,
            in1 => \N__15765\,
            in2 => \N__19736\,
            in3 => \N__15405\,
            lcout => \Lab_UT.dictrl.g0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__19714\,
            in1 => \N__19112\,
            in2 => \N__19921\,
            in3 => \N__19779\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_x1_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19454\,
            in1 => \N__20007\,
            in2 => \N__15784\,
            in3 => \N__15710\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m22_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_ns_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15415\,
            in3 => \N__15248\,
            lcout => \Lab_UT.dictrl.N_72_mux\,
            ltout => \Lab_UT.dictrl.N_72_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19868\,
            in2 => \N__15412\,
            in3 => \N__19778\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__15795\,
            in1 => \N__19464\,
            in2 => \N__19545\,
            in3 => \N__15409\,
            lcout => \Lab_UT.dictrl.g0_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_x1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19513\,
            in1 => \N__15621\,
            in2 => \N__15331\,
            in3 => \N__15299\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15280\,
            in3 => \N__15277\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15232\,
            in1 => \N__15268\,
            in2 => \N__15262\,
            in3 => \N__21426\,
            lcout => \Lab_UT.dictrl.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15647\,
            in1 => \N__19398\,
            in2 => \N__15625\,
            in3 => \N__19363\,
            lcout => \Lab_UT.dictrl.m22Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__19364\,
            in1 => \N__15623\,
            in2 => \N__19405\,
            in3 => \N__19691\,
            lcout => \Lab_UT.dictrl.g0_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20032\,
            in1 => \N__21431\,
            in2 => \N__15799\,
            in3 => \N__15709\,
            lcout => \G_6_0_a6_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19399\,
            in1 => \N__15622\,
            in2 => \N__19544\,
            in3 => \N__15648\,
            lcout => \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_rep1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15601\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__15474\,
            sr => \N__20973\
        );

    \buart.Z_rx.shifter_7_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15600\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__15474\,
            sr => \N__20973\
        );

    \buart.Z_rx.shifter_fast_0_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20191\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__15474\,
            sr => \N__20973\
        );

    \buart.Z_rx.shifter_6_rep1_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15525\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => \N__15474\,
            sr => \N__20973\
        );

    \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15988\,
            in1 => \N__20739\,
            in2 => \N__15448\,
            in3 => \N__15967\,
            lcout => \uu2.un3_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__15969\,
            in1 => \N__15993\,
            in2 => \N__21952\,
            in3 => \N__20741\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15853\,
            sr => \N__15841\
        );

    \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16012\,
            in1 => \N__15866\,
            in2 => \_gnd_net_\,
            in3 => \N__21946\,
            lcout => OPEN,
            ltout => \uu2.un3_w_addr_user_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIINVH_4_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16048\,
            in1 => \N__16189\,
            in2 => \N__16162\,
            in3 => \N__16159\,
            lcout => \uu2.un3_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15989\,
            in1 => \N__21903\,
            in2 => \_gnd_net_\,
            in3 => \N__16137\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_7_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__16049\,
            in1 => \N__15915\,
            in2 => \N__16018\,
            in3 => \N__15903\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15853\,
            sr => \N__15841\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20740\,
            in1 => \N__21947\,
            in2 => \N__15994\,
            in3 => \N__15968\,
            lcout => \uu2.un404_ci\,
            ltout => \uu2.un404_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__15867\,
            in1 => \N__15902\,
            in2 => \N__15880\,
            in3 => \N__15877\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__15853\,
            sr => \N__15841\
        );

    \uu2.bitmap_290_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100111"
        )
    port map (
            in0 => \N__16557\,
            in1 => \N__16379\,
            in2 => \N__17372\,
            in3 => \N__16416\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_194_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__16415\,
            in1 => \N__17359\,
            in2 => \N__16388\,
            in3 => \N__16556\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_66_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000110101"
        )
    port map (
            in0 => \N__16559\,
            in1 => \N__16383\,
            in2 => \N__17373\,
            in3 => \N__16418\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_RNIPDM31_66_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__15811\,
            in1 => \N__16309\,
            in2 => \N__16264\,
            in3 => \N__15805\,
            lcout => \uu2.bitmap_pmux_20_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000110110"
        )
    port map (
            in0 => \N__16555\,
            in1 => \N__16375\,
            in2 => \N__17371\,
            in3 => \N__16414\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_34_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111101111001"
        )
    port map (
            in0 => \N__16417\,
            in1 => \N__17363\,
            in2 => \N__16389\,
            in3 => \N__16558\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_RNIP2JO1_34_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001010"
        )
    port map (
            in0 => \N__16492\,
            in1 => \N__16486\,
            in2 => \N__16480\,
            in3 => \N__16463\,
            lcout => \uu2.bitmap_RNIP2JO1Z0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_69_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__16419\,
            in1 => \N__17367\,
            in2 => \N__16390\,
            in3 => \N__16560\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__20906\
        );

    \uu2.bitmap_314_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011101"
        )
    port map (
            in0 => \N__16803\,
            in1 => \N__16840\,
            in2 => \N__16883\,
            in3 => \N__16908\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20904\
        );

    \uu2.bitmap_218_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010101"
        )
    port map (
            in0 => \N__16907\,
            in1 => \N__16870\,
            in2 => \N__16845\,
            in3 => \N__16802\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20904\
        );

    \uu2.bitmap_90_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__16805\,
            in1 => \N__16844\,
            in2 => \N__16884\,
            in3 => \N__16910\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20904\
        );

    \uu2.bitmap_RNIJ4K41_90_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__16310\,
            in1 => \N__16270\,
            in2 => \N__16250\,
            in3 => \N__16204\,
            lcout => \uu2.bitmap_pmux_19_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__16801\,
            in1 => \N__16836\,
            in2 => \N__16882\,
            in3 => \N__16906\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20904\
        );

    \uu2.bitmap_58_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__16909\,
            in1 => \N__16874\,
            in2 => \N__16846\,
            in3 => \N__16804\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__20904\
        );

    \uu2.bitmap_RNIM5E21_314_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16779\,
            in1 => \N__16765\,
            in2 => \_gnd_net_\,
            in3 => \N__16681\,
            lcout => \uu2.bitmap_RNIM5E21Z0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIKGSI_58_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16713\,
            in1 => \N__16693\,
            in2 => \_gnd_net_\,
            in3 => \N__16687\,
            lcout => \uu2.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__17968\,
            in1 => \N__17530\,
            in2 => \N__18011\,
            in3 => \N__17176\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI62AM_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16675\,
            in2 => \_gnd_net_\,
            in3 => \N__17869\,
            lcout => \Lab_UT.didp.un1_dicLdStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17518\,
            in1 => \N__16624\,
            in2 => \_gnd_net_\,
            in3 => \N__16591\,
            lcout => \Lab_UT.min1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17108\,
            in1 => \N__20341\,
            in2 => \N__16528\,
            in3 => \N__17433\,
            lcout => \Lab_UT.didp.countrce4.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17002\,
            in1 => \N__17231\,
            in2 => \_gnd_net_\,
            in3 => \N__17933\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__16941\,
            in1 => \N__20524\,
            in2 => \N__17533\,
            in3 => \N__17175\,
            lcout => \Lab_UT.didp.countrce3.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17727\,
            in2 => \_gnd_net_\,
            in3 => \N__17582\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17639\,
            in1 => \N__20340\,
            in2 => \N__17524\,
            in3 => \N__17269\,
            lcout => \Lab_UT.didp.countrce1.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17499\,
            in1 => \N__17430\,
            in2 => \_gnd_net_\,
            in3 => \N__17401\,
            lcout => \Lab_UT.min1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__17746\,
            in1 => \N__17329\,
            in2 => \N__17323\,
            in3 => \N__17270\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17000\,
            in1 => \N__17236\,
            in2 => \N__17187\,
            in3 => \N__17930\,
            lcout => \Lab_UT.didp.countrce3.ce_12_0_a6_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17117\,
            in1 => \N__20516\,
            in2 => \N__17059\,
            in3 => \N__17040\,
            lcout => \Lab_UT.didp.countrce4.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__20200\,
            in2 => \N__16953\,
            in3 => \N__17931\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17932\,
            in1 => \N__18012\,
            in2 => \N__17971\,
            in3 => \N__17964\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_esr_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18169\,
            in1 => \N__17827\,
            in2 => \N__18861\,
            in3 => \N__18120\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__18526\,
            sr => \N__20946\
        );

    \Lab_UT.dictrl.state_ret_11_ess_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__18121\,
            in1 => \N__18857\,
            in2 => \N__17835\,
            in3 => \N__18170\,
            lcout => \Lab_UT.LdSones_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__18526\,
            sr => \N__20946\
        );

    \Lab_UT.dictrl.state_ret_8_ess_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__18171\,
            in1 => \N__17831\,
            in2 => \N__18862\,
            in3 => \N__18122\,
            lcout => \Lab_UT.state_ret_8_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__18526\,
            sr => \N__20946\
        );

    \Lab_UT.didp.state_ret_1_esr_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__18123\,
            in1 => \_gnd_net_\,
            in2 => \N__17836\,
            in3 => \N__18172\,
            lcout => \Lab_UT.didp.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__18526\,
            sr => \N__20946\
        );

    \Lab_UT.didp.ce_RNIFQ9K_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__17779\,
            in1 => \N__17770\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.un1_dicLdSones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__17726\,
            in1 => \N__20186\,
            in2 => \N__17638\,
            in3 => \N__17589\,
            lcout => \Lab_UT.didp.countrce1.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__18495\,
            in1 => \N__21486\,
            in2 => \_gnd_net_\,
            in3 => \N__18670\,
            lcout => \Lab_UT.next_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI81O17_2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__19259\,
            in1 => \N__21307\,
            in2 => \N__18597\,
            in3 => \N__21229\,
            lcout => \Lab_UT.dictrl.g0_1_mb_rn_0\,
            ltout => \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__18496\,
            in1 => \_gnd_net_\,
            in2 => \N__18664\,
            in3 => \N__21487\,
            lcout => \Lab_UT.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22306\,
            ce => \N__18537\,
            sr => \N__20940\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__21108\,
            in1 => \N__18657\,
            in2 => \N__18630\,
            in3 => \N__21230\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18593\,
            in2 => \N__18565\,
            in3 => \N__19263\,
            lcout => \Lab_UT.dictrl.state_i_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22306\,
            ce => \N__18537\,
            sr => \N__20940\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__21107\,
            in1 => \_gnd_net_\,
            in2 => \N__19274\,
            in3 => \N__21228\,
            lcout => \Lab_UT.dictrl.g0_1_mb_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18482\,
            in2 => \_gnd_net_\,
            in3 => \N__21106\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un15_loadalarm_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__18920\,
            in1 => \N__21227\,
            in2 => \N__18466\,
            in3 => \N__20583\,
            lcout => \Lab_UT.dictrl.loadalarm_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18457\,
            in1 => \N__18216\,
            in2 => \_gnd_net_\,
            in3 => \N__18370\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22297\,
            ce => 'H',
            sr => \N__20947\
        );

    \Lab_UT.dictrl.state_ret_9_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__18153\,
            in1 => \N__18118\,
            in2 => \N__18088\,
            in3 => \N__18935\,
            lcout => \Lab_UT.dicLdSones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22297\,
            ce => 'H',
            sr => \N__20947\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21250\,
            in2 => \_gnd_net_\,
            in3 => \N__21373\,
            lcout => \Lab_UT.dictrl.m34_0\,
            ltout => \Lab_UT.dictrl.m34_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m35_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__18801\,
            in1 => \N__18777\,
            in2 => \N__18889\,
            in3 => \N__21141\,
            lcout => \Lab_UT.dictrl.next_state_1_3\,
            ltout => \Lab_UT.dictrl.next_state_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18726\,
            in2 => \N__18865\,
            in3 => \N__19231\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19229\,
            in1 => \N__19030\,
            in2 => \_gnd_net_\,
            in3 => \N__21139\,
            lcout => \Lab_UT.dictrl.N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21140\,
            in1 => \N__19230\,
            in2 => \_gnd_net_\,
            in3 => \N__19034\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__21374\,
            in1 => \N__18829\,
            in2 => \N__18820\,
            in3 => \N__19555\,
            lcout => \Lab_UT.dictrl.N_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21142\,
            in1 => \N__18802\,
            in2 => \N__18787\,
            in3 => \N__18778\,
            lcout => \Lab_UT.dictrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22289\,
            ce => \N__19327\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__20532\,
            in1 => \_gnd_net_\,
            in2 => \N__18970\,
            in3 => \N__21418\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18695\,
            in2 => \N__19345\,
            in3 => \N__18895\,
            lcout => \Lab_UT.dictrl.next_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => \N__19341\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__19290\,
            in1 => \N__19264\,
            in2 => \_gnd_net_\,
            in3 => \N__21417\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_latmux_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__19265\,
            in1 => \N__18965\,
            in2 => \N__19141\,
            in3 => \N__20533\,
            lcout => \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m7_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19123\,
            in2 => \_gnd_net_\,
            in3 => \N__19826\,
            lcout => \Lab_UT.dictrl.N_8_0\,
            ltout => \Lab_UT.dictrl.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__20498\,
            in1 => \N__20352\,
            in2 => \N__19096\,
            in3 => \N__20618\,
            lcout => \Lab_UT.dictrl.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101110000"
        )
    port map (
            in0 => \N__20617\,
            in1 => \N__18937\,
            in2 => \N__19072\,
            in3 => \N__21416\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_6_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000000100"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__19068\,
            in2 => \N__19093\,
            in3 => \N__19930\,
            lcout => \Lab_UT.dictrl.G_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__19084\,
            in1 => \N__19078\,
            in2 => \N__20517\,
            in3 => \N__20620\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.i8_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000101"
        )
    port map (
            in0 => \N__19069\,
            in1 => \N__18969\,
            in2 => \N__18952\,
            in3 => \N__18938\,
            lcout => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__20358\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__20619\,
            lcout => \Lab_UT.dictrl.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m14_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__19824\,
            in1 => \N__20494\,
            in2 => \_gnd_net_\,
            in3 => \N__19597\,
            lcout => \Lab_UT.dictrl.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__20302\,
            in1 => \N__19825\,
            in2 => \N__20198\,
            in3 => \N__20031\,
            lcout => \G_6_0_a6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__19918\,
            in1 => \N__19823\,
            in2 => \N__19737\,
            in3 => \N__19627\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19606\,
            in2 => \N__19600\,
            in3 => \N__19596\,
            lcout => \Lab_UT.dictrl.N_59_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19546\,
            in1 => \N__19512\,
            in2 => \_gnd_net_\,
            in3 => \N__19498\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__19477\,
            in1 => \N__19465\,
            in2 => \N__19408\,
            in3 => \N__19404\,
            lcout => \Lab_UT.dictrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19372\,
            lcout => \Lab_UT.dictrl.g0_6_3\,
            ltout => \Lab_UT.dictrl.g0_6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__21456\,
            in1 => \N__21466\,
            in2 => \N__21490\,
            in3 => \N__21442\,
            lcout => \Lab_UT.dictrl.N_57_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_8_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__21472\,
            in1 => \N__21465\,
            in2 => \N__21457\,
            in3 => \N__21441\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_13_RNO_4_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101110111"
        )
    port map (
            in0 => \N__21303\,
            in1 => \N__21283\,
            in2 => \N__21172\,
            in3 => \N__21153\,
            lcout => \Lab_UT.dictrl.G_25_i_a5_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111111100"
        )
    port map (
            in0 => \N__21517\,
            in1 => \N__21556\,
            in2 => \N__21714\,
            in3 => \N__21578\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \N__20974\
        );

    \buart.Z_tx.bitcount_0_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21577\,
            in1 => \N__21698\,
            in2 => \_gnd_net_\,
            in3 => \N__21516\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \N__20974\
        );

    \buart.Z_tx.bitcount_3_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__21595\,
            in1 => \N__21496\,
            in2 => \N__21715\,
            in3 => \N__21580\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \N__20974\
        );

    \buart.Z_tx.bitcount_2_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010110"
        )
    port map (
            in0 => \N__21579\,
            in1 => \N__21721\,
            in2 => \N__21538\,
            in3 => \N__21702\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \N__20974\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20742\,
            in1 => \N__21917\,
            in2 => \_gnd_net_\,
            in3 => \N__20704\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21951\,
            in1 => \N__21918\,
            in2 => \_gnd_net_\,
            in3 => \N__21799\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__21514\,
            in1 => \N__21554\,
            in2 => \_gnd_net_\,
            in3 => \N__21575\,
            lcout => \buart.Z_tx.un1_bitcount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22027\,
            in2 => \_gnd_net_\,
            in3 => \N__22011\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21678\,
            in2 => \_gnd_net_\,
            in3 => \N__21576\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22010\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21594\,
            in2 => \_gnd_net_\,
            in3 => \N__21513\,
            lcout => OPEN,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__21533\,
            in1 => \N__21553\,
            in2 => \N__21583\,
            in3 => \N__21967\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__21555\,
            in1 => \N__21534\,
            in2 => \N__21520\,
            in3 => \N__21515\,
            lcout => \buart.Z_tx.un1_bitcount_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22026\,
            in2 => \N__22012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21991\,
            in3 => \N__22372\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__22350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21969\,
            in1 => \N__22036\,
            in2 => \_gnd_net_\,
            in3 => \N__22369\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__22350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22063\,
            in3 => \N__22366\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__22350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__21970\,
            in1 => \_gnd_net_\,
            in2 => \N__22075\,
            in3 => \N__22363\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__22350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__22050\,
            in1 => \N__21968\,
            in2 => \_gnd_net_\,
            in3 => \N__22360\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__22071\,
            in1 => \N__22059\,
            in2 => \N__22051\,
            in3 => \N__22035\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22025\,
            in1 => \N__22006\,
            in2 => \N__21990\,
            in3 => \N__21976\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
