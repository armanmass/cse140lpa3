// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 21 2019 00:12:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__22472;
    wire N__22471;
    wire N__22470;
    wire N__22463;
    wire N__22462;
    wire N__22461;
    wire N__22454;
    wire N__22453;
    wire N__22452;
    wire N__22445;
    wire N__22444;
    wire N__22443;
    wire N__22436;
    wire N__22435;
    wire N__22434;
    wire N__22427;
    wire N__22426;
    wire N__22425;
    wire N__22418;
    wire N__22417;
    wire N__22416;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22400;
    wire N__22399;
    wire N__22398;
    wire N__22391;
    wire N__22390;
    wire N__22389;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22350;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22346;
    wire N__22345;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22337;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22330;
    wire N__22329;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22317;
    wire N__22316;
    wire N__22315;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22311;
    wire N__22310;
    wire N__22309;
    wire N__22308;
    wire N__22307;
    wire N__22306;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22301;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22275;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22260;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22071;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22054;
    wire N__22051;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22036;
    wire N__22035;
    wire N__22030;
    wire N__22027;
    wire N__22026;
    wire N__22025;
    wire N__22022;
    wire N__22017;
    wire N__22012;
    wire N__22011;
    wire N__22010;
    wire N__22007;
    wire N__22006;
    wire N__22001;
    wire N__21996;
    wire N__21991;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21969;
    wire N__21968;
    wire N__21967;
    wire N__21960;
    wire N__21957;
    wire N__21952;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21942;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21911;
    wire N__21910;
    wire N__21909;
    wire N__21904;
    wire N__21903;
    wire N__21902;
    wire N__21901;
    wire N__21900;
    wire N__21899;
    wire N__21886;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21874;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21784;
    wire N__21783;
    wire N__21782;
    wire N__21781;
    wire N__21780;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21773;
    wire N__21770;
    wire N__21761;
    wire N__21756;
    wire N__21753;
    wire N__21744;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21707;
    wire N__21706;
    wire N__21703;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21679;
    wire N__21678;
    wire N__21669;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21631;
    wire N__21622;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21595;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21583;
    wire N__21580;
    wire N__21579;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21566;
    wire N__21561;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21553;
    wire N__21550;
    wire N__21543;
    wire N__21538;
    wire N__21535;
    wire N__21534;
    wire N__21533;
    wire N__21530;
    wire N__21525;
    wire N__21520;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21508;
    wire N__21501;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21486;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21465;
    wire N__21460;
    wire N__21457;
    wire N__21456;
    wire N__21453;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21419;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21382;
    wire N__21377;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21373;
    wire N__21368;
    wire N__21365;
    wire N__21360;
    wire N__21359;
    wire N__21344;
    wire N__21339;
    wire N__21334;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21318;
    wire N__21307;
    wire N__21304;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21289;
    wire N__21288;
    wire N__21287;
    wire N__21284;
    wire N__21283;
    wire N__21282;
    wire N__21279;
    wire N__21278;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21236;
    wire N__21231;
    wire N__21230;
    wire N__21229;
    wire N__21228;
    wire N__21227;
    wire N__21226;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21211;
    wire N__21204;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21172;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21165;
    wire N__21160;
    wire N__21159;
    wire N__21154;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21136;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21092;
    wire N__21085;
    wire N__21080;
    wire N__21073;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21025;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20994;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20973;
    wire N__20972;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20965;
    wire N__20964;
    wire N__20963;
    wire N__20962;
    wire N__20961;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20955;
    wire N__20954;
    wire N__20953;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20906;
    wire N__20905;
    wire N__20904;
    wire N__20903;
    wire N__20902;
    wire N__20901;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20897;
    wire N__20896;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20742;
    wire N__20741;
    wire N__20740;
    wire N__20739;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20727;
    wire N__20724;
    wire N__20719;
    wire N__20716;
    wire N__20711;
    wire N__20704;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20674;
    wire N__20663;
    wire N__20660;
    wire N__20653;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20623;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20618;
    wire N__20617;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20599;
    wire N__20596;
    wire N__20587;
    wire N__20584;
    wire N__20583;
    wire N__20582;
    wire N__20579;
    wire N__20574;
    wire N__20569;
    wire N__20566;
    wire N__20561;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20533;
    wire N__20532;
    wire N__20527;
    wire N__20524;
    wire N__20523;
    wire N__20522;
    wire N__20521;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20512;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20498;
    wire N__20495;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20483;
    wire N__20478;
    wire N__20475;
    wire N__20470;
    wire N__20469;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20461;
    wire N__20460;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20442;
    wire N__20441;
    wire N__20438;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20419;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20400;
    wire N__20397;
    wire N__20392;
    wire N__20383;
    wire N__20380;
    wire N__20359;
    wire N__20358;
    wire N__20353;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20341;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20331;
    wire N__20330;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20312;
    wire N__20311;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20303;
    wire N__20302;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20287;
    wire N__20284;
    wire N__20279;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20262;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20248;
    wire N__20241;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20220;
    wire N__20213;
    wire N__20200;
    wire N__20199;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20191;
    wire N__20188;
    wire N__20187;
    wire N__20186;
    wire N__20185;
    wire N__20184;
    wire N__20183;
    wire N__20178;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20127;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20110;
    wire N__20107;
    wire N__20100;
    wire N__20091;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20053;
    wire N__20038;
    wire N__20037;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20030;
    wire N__20029;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20015;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19991;
    wire N__19990;
    wire N__19987;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19969;
    wire N__19966;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19946;
    wire N__19943;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19920;
    wire N__19919;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19908;
    wire N__19907;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19895;
    wire N__19894;
    wire N__19891;
    wire N__19886;
    wire N__19881;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19869;
    wire N__19868;
    wire N__19865;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19835;
    wire N__19828;
    wire N__19827;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19811;
    wire N__19808;
    wire N__19801;
    wire N__19800;
    wire N__19795;
    wire N__19790;
    wire N__19783;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19762;
    wire N__19759;
    wire N__19754;
    wire N__19751;
    wire N__19738;
    wire N__19737;
    wire N__19736;
    wire N__19735;
    wire N__19732;
    wire N__19731;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19720;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19656;
    wire N__19653;
    wire N__19646;
    wire N__19643;
    wire N__19636;
    wire N__19633;
    wire N__19632;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19596;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19579;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19518;
    wire N__19513;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19498;
    wire N__19495;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19454;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19446;
    wire N__19443;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19420;
    wire N__19417;
    wire N__19408;
    wire N__19405;
    wire N__19404;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19385;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19352;
    wire N__19345;
    wire N__19342;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19331;
    wire N__19328;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19294;
    wire N__19291;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19276;
    wire N__19275;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19266;
    wire N__19265;
    wire N__19264;
    wire N__19263;
    wire N__19260;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19239;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19192;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19176;
    wire N__19173;
    wire N__19168;
    wire N__19161;
    wire N__19158;
    wire N__19141;
    wire N__19138;
    wire N__19137;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19122;
    wire N__19121;
    wire N__19118;
    wire N__19113;
    wire N__19112;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19069;
    wire N__19068;
    wire N__19065;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19052;
    wire N__19051;
    wire N__19050;
    wire N__19049;
    wire N__19042;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19008;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18989;
    wire N__18970;
    wire N__18969;
    wire N__18966;
    wire N__18965;
    wire N__18962;
    wire N__18957;
    wire N__18952;
    wire N__18949;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18907;
    wire N__18904;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18879;
    wire N__18878;
    wire N__18875;
    wire N__18870;
    wire N__18865;
    wire N__18862;
    wire N__18861;
    wire N__18858;
    wire N__18857;
    wire N__18854;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18840;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18816;
    wire N__18815;
    wire N__18814;
    wire N__18805;
    wire N__18802;
    wire N__18801;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18770;
    wire N__18769;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18750;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18726;
    wire N__18723;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18700;
    wire N__18699;
    wire N__18696;
    wire N__18695;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18634;
    wire N__18631;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18597;
    wire N__18594;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18565;
    wire N__18562;
    wire N__18561;
    wire N__18560;
    wire N__18559;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18538;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18530;
    wire N__18527;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18509;
    wire N__18506;
    wire N__18501;
    wire N__18496;
    wire N__18495;
    wire N__18490;
    wire N__18487;
    wire N__18486;
    wire N__18483;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18456;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18448;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18426;
    wire N__18423;
    wire N__18418;
    wire N__18417;
    wire N__18416;
    wire N__18415;
    wire N__18412;
    wire N__18405;
    wire N__18402;
    wire N__18395;
    wire N__18390;
    wire N__18383;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18365;
    wire N__18364;
    wire N__18363;
    wire N__18362;
    wire N__18361;
    wire N__18360;
    wire N__18359;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18351;
    wire N__18350;
    wire N__18349;
    wire N__18346;
    wire N__18341;
    wire N__18332;
    wire N__18327;
    wire N__18326;
    wire N__18325;
    wire N__18324;
    wire N__18321;
    wire N__18320;
    wire N__18319;
    wire N__18316;
    wire N__18311;
    wire N__18308;
    wire N__18301;
    wire N__18294;
    wire N__18291;
    wire N__18286;
    wire N__18283;
    wire N__18268;
    wire N__18267;
    wire N__18266;
    wire N__18265;
    wire N__18262;
    wire N__18261;
    wire N__18260;
    wire N__18253;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18244;
    wire N__18243;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18222;
    wire N__18217;
    wire N__18216;
    wire N__18213;
    wire N__18208;
    wire N__18203;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18172;
    wire N__18171;
    wire N__18170;
    wire N__18169;
    wire N__18160;
    wire N__18159;
    wire N__18158;
    wire N__18157;
    wire N__18154;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18133;
    wire N__18124;
    wire N__18123;
    wire N__18122;
    wire N__18121;
    wire N__18120;
    wire N__18119;
    wire N__18118;
    wire N__18115;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18088;
    wire N__18087;
    wire N__18084;
    wire N__18083;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18075;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18062;
    wire N__18057;
    wire N__18050;
    wire N__18047;
    wire N__18046;
    wire N__18041;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18023;
    wire N__18020;
    wire N__18013;
    wire N__18012;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17989;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17941;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17933;
    wire N__17932;
    wire N__17931;
    wire N__17930;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17913;
    wire N__17910;
    wire N__17905;
    wire N__17896;
    wire N__17895;
    wire N__17894;
    wire N__17891;
    wire N__17890;
    wire N__17889;
    wire N__17886;
    wire N__17881;
    wire N__17878;
    wire N__17873;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17843;
    wire N__17836;
    wire N__17835;
    wire N__17832;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17826;
    wire N__17825;
    wire N__17824;
    wire N__17815;
    wire N__17810;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17728;
    wire N__17727;
    wire N__17726;
    wire N__17725;
    wire N__17722;
    wire N__17721;
    wire N__17718;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17689;
    wire N__17688;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17667;
    wire N__17664;
    wire N__17659;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17639;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17605;
    wire N__17604;
    wire N__17603;
    wire N__17602;
    wire N__17595;
    wire N__17592;
    wire N__17591;
    wire N__17590;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17582;
    wire N__17579;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17520;
    wire N__17519;
    wire N__17518;
    wire N__17511;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17505;
    wire N__17504;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17479;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17456;
    wire N__17451;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17433;
    wire N__17432;
    wire N__17431;
    wire N__17430;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17401;
    wire N__17398;
    wire N__17397;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17374;
    wire N__17373;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17367;
    wire N__17364;
    wire N__17363;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17302;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17286;
    wire N__17283;
    wire N__17278;
    wire N__17277;
    wire N__17272;
    wire N__17271;
    wire N__17270;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17236;
    wire N__17235;
    wire N__17232;
    wire N__17231;
    wire N__17228;
    wire N__17227;
    wire N__17226;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17197;
    wire N__17188;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17143;
    wire N__17142;
    wire N__17141;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17121;
    wire N__17118;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17110;
    wire N__17109;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17046;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16997;
    wire N__16996;
    wire N__16995;
    wire N__16994;
    wire N__16989;
    wire N__16986;
    wire N__16985;
    wire N__16982;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16957;
    wire N__16956;
    wire N__16955;
    wire N__16954;
    wire N__16953;
    wire N__16950;
    wire N__16945;
    wire N__16942;
    wire N__16941;
    wire N__16938;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16912;
    wire N__16911;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16901;
    wire N__16890;
    wire N__16885;
    wire N__16884;
    wire N__16883;
    wire N__16882;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16874;
    wire N__16871;
    wire N__16870;
    wire N__16867;
    wire N__16862;
    wire N__16851;
    wire N__16846;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16836;
    wire N__16835;
    wire N__16834;
    wire N__16823;
    wire N__16818;
    wire N__16815;
    wire N__16810;
    wire N__16807;
    wire N__16806;
    wire N__16805;
    wire N__16804;
    wire N__16803;
    wire N__16802;
    wire N__16801;
    wire N__16796;
    wire N__16785;
    wire N__16780;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16765;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16739;
    wire N__16732;
    wire N__16731;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16714;
    wire N__16713;
    wire N__16710;
    wire N__16703;
    wire N__16700;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16657;
    wire N__16656;
    wire N__16651;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16639;
    wire N__16636;
    wire N__16635;
    wire N__16634;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16624;
    wire N__16621;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16591;
    wire N__16590;
    wire N__16587;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16569;
    wire N__16564;
    wire N__16561;
    wire N__16560;
    wire N__16559;
    wire N__16558;
    wire N__16557;
    wire N__16556;
    wire N__16555;
    wire N__16552;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16467;
    wire N__16464;
    wire N__16463;
    wire N__16462;
    wire N__16459;
    wire N__16458;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16446;
    wire N__16441;
    wire N__16436;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16419;
    wire N__16418;
    wire N__16417;
    wire N__16416;
    wire N__16415;
    wire N__16414;
    wire N__16411;
    wire N__16398;
    wire N__16395;
    wire N__16390;
    wire N__16389;
    wire N__16388;
    wire N__16387;
    wire N__16384;
    wire N__16383;
    wire N__16380;
    wire N__16379;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16332;
    wire N__16331;
    wire N__16326;
    wire N__16325;
    wire N__16324;
    wire N__16323;
    wire N__16322;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16299;
    wire N__16294;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16263;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16251;
    wire N__16250;
    wire N__16249;
    wire N__16246;
    wire N__16237;
    wire N__16236;
    wire N__16235;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16223;
    wire N__16216;
    wire N__16213;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16188;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16182;
    wire N__16177;
    wire N__16172;
    wire N__16167;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16152;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16137;
    wire N__16136;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16128;
    wire N__16127;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16112;
    wire N__16111;
    wire N__16108;
    wire N__16103;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16084;
    wire N__16081;
    wire N__16072;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16036;
    wire N__16033;
    wire N__16026;
    wire N__16023;
    wire N__16018;
    wire N__16015;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16009;
    wire N__16004;
    wire N__16001;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15969;
    wire N__15968;
    wire N__15967;
    wire N__15966;
    wire N__15963;
    wire N__15962;
    wire N__15961;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15943;
    wire N__15940;
    wire N__15935;
    wire N__15928;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15916;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15899;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15867;
    wire N__15866;
    wire N__15863;
    wire N__15858;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15823;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15811;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15795;
    wire N__15790;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15786;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15780;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15727;
    wire N__15724;
    wire N__15715;
    wire N__15712;
    wire N__15711;
    wire N__15710;
    wire N__15709;
    wire N__15708;
    wire N__15705;
    wire N__15700;
    wire N__15699;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15687;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15648;
    wire N__15647;
    wire N__15646;
    wire N__15645;
    wire N__15642;
    wire N__15637;
    wire N__15632;
    wire N__15625;
    wire N__15624;
    wire N__15623;
    wire N__15622;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15606;
    wire N__15601;
    wire N__15600;
    wire N__15599;
    wire N__15594;
    wire N__15591;
    wire N__15586;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15568;
    wire N__15565;
    wire N__15564;
    wire N__15563;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15554;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15536;
    wire N__15533;
    wire N__15526;
    wire N__15525;
    wire N__15524;
    wire N__15521;
    wire N__15512;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15481;
    wire N__15480;
    wire N__15479;
    wire N__15478;
    wire N__15477;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15444;
    wire N__15443;
    wire N__15440;
    wire N__15439;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15405;
    wire N__15404;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15389;
    wire N__15388;
    wire N__15387;
    wire N__15386;
    wire N__15385;
    wire N__15384;
    wire N__15379;
    wire N__15378;
    wire N__15377;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15361;
    wire N__15354;
    wire N__15351;
    wire N__15346;
    wire N__15331;
    wire N__15328;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15307;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15299;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15258;
    wire N__15257;
    wire N__15252;
    wire N__15249;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15225;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15215;
    wire N__15212;
    wire N__15207;
    wire N__15202;
    wire N__15199;
    wire N__15198;
    wire N__15195;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15186;
    wire N__15185;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15169;
    wire N__15162;
    wire N__15159;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15047;
    wire N__15046;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14982;
    wire N__14977;
    wire N__14974;
    wire N__14973;
    wire N__14972;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14904;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14892;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14871;
    wire N__14868;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14848;
    wire N__14845;
    wire N__14844;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14809;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14773;
    wire N__14772;
    wire N__14771;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14747;
    wire N__14746;
    wire N__14743;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14721;
    wire N__14718;
    wire N__14713;
    wire N__14712;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14667;
    wire N__14666;
    wire N__14659;
    wire N__14658;
    wire N__14657;
    wire N__14654;
    wire N__14649;
    wire N__14648;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14636;
    wire N__14629;
    wire N__14628;
    wire N__14627;
    wire N__14626;
    wire N__14623;
    wire N__14622;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14610;
    wire N__14609;
    wire N__14606;
    wire N__14599;
    wire N__14596;
    wire N__14591;
    wire N__14584;
    wire N__14583;
    wire N__14578;
    wire N__14577;
    wire N__14576;
    wire N__14575;
    wire N__14572;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14552;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14506;
    wire N__14503;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14499;
    wire N__14492;
    wire N__14489;
    wire N__14488;
    wire N__14485;
    wire N__14484;
    wire N__14481;
    wire N__14476;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14455;
    wire N__14452;
    wire N__14451;
    wire N__14450;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14438;
    wire N__14437;
    wire N__14434;
    wire N__14433;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14415;
    wire N__14412;
    wire N__14401;
    wire N__14400;
    wire N__14397;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14379;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14358;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14347;
    wire N__14344;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14326;
    wire N__14323;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14301;
    wire N__14300;
    wire N__14299;
    wire N__14298;
    wire N__14297;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14285;
    wire N__14278;
    wire N__14275;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14258;
    wire N__14257;
    wire N__14254;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14224;
    wire N__14223;
    wire N__14222;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14216;
    wire N__14211;
    wire N__14206;
    wire N__14201;
    wire N__14196;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14178;
    wire N__14173;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14154;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14139;
    wire N__14134;
    wire N__14133;
    wire N__14132;
    wire N__14131;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14117;
    wire N__14116;
    wire N__14113;
    wire N__14100;
    wire N__14095;
    wire N__14094;
    wire N__14093;
    wire N__14092;
    wire N__14091;
    wire N__14090;
    wire N__14089;
    wire N__14086;
    wire N__14073;
    wire N__14068;
    wire N__14067;
    wire N__14066;
    wire N__14065;
    wire N__14064;
    wire N__14063;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14029;
    wire N__14028;
    wire N__14027;
    wire N__14026;
    wire N__14025;
    wire N__14024;
    wire N__14023;
    wire N__14020;
    wire N__14007;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13983;
    wire N__13982;
    wire N__13979;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13959;
    wire N__13958;
    wire N__13957;
    wire N__13954;
    wire N__13953;
    wire N__13948;
    wire N__13947;
    wire N__13946;
    wire N__13945;
    wire N__13944;
    wire N__13943;
    wire N__13936;
    wire N__13933;
    wire N__13932;
    wire N__13925;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13900;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13827;
    wire N__13826;
    wire N__13823;
    wire N__13818;
    wire N__13813;
    wire N__13810;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13785;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13765;
    wire N__13764;
    wire N__13761;
    wire N__13760;
    wire N__13759;
    wire N__13758;
    wire N__13757;
    wire N__13754;
    wire N__13753;
    wire N__13752;
    wire N__13751;
    wire N__13750;
    wire N__13749;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13721;
    wire N__13716;
    wire N__13713;
    wire N__13706;
    wire N__13703;
    wire N__13698;
    wire N__13691;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13662;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13639;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13614;
    wire N__13609;
    wire N__13608;
    wire N__13607;
    wire N__13606;
    wire N__13603;
    wire N__13602;
    wire N__13601;
    wire N__13596;
    wire N__13595;
    wire N__13590;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13563;
    wire N__13560;
    wire N__13559;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13547;
    wire N__13546;
    wire N__13543;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13498;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13470;
    wire N__13469;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13463;
    wire N__13462;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13438;
    wire N__13435;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13393;
    wire N__13392;
    wire N__13391;
    wire N__13388;
    wire N__13383;
    wire N__13380;
    wire N__13375;
    wire N__13372;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13342;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13338;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13326;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13312;
    wire N__13311;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13283;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13233;
    wire N__13228;
    wire N__13225;
    wire N__13224;
    wire N__13221;
    wire N__13220;
    wire N__13219;
    wire N__13216;
    wire N__13215;
    wire N__13214;
    wire N__13211;
    wire N__13204;
    wire N__13199;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13176;
    wire N__13175;
    wire N__13174;
    wire N__13173;
    wire N__13172;
    wire N__13171;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13152;
    wire N__13147;
    wire N__13142;
    wire N__13139;
    wire N__13134;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13096;
    wire N__13091;
    wire N__13082;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13051;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13028;
    wire N__13025;
    wire N__13024;
    wire N__13023;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13008;
    wire N__13005;
    wire N__12994;
    wire N__12993;
    wire N__12992;
    wire N__12991;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12964;
    wire N__12963;
    wire N__12962;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12956;
    wire N__12953;
    wire N__12952;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12938;
    wire N__12937;
    wire N__12934;
    wire N__12933;
    wire N__12930;
    wire N__12925;
    wire N__12920;
    wire N__12913;
    wire N__12906;
    wire N__12895;
    wire N__12894;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12886;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12880;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12868;
    wire N__12867;
    wire N__12866;
    wire N__12865;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12851;
    wire N__12844;
    wire N__12837;
    wire N__12826;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12805;
    wire N__12804;
    wire N__12797;
    wire N__12796;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12780;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12741;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12729;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12683;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12603;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12512;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12465;
    wire N__12460;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12442;
    wire N__12439;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12395;
    wire N__12394;
    wire N__12391;
    wire N__12384;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12369;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12354;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12285;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12256;
    wire N__12255;
    wire N__12254;
    wire N__12253;
    wire N__12252;
    wire N__12249;
    wire N__12248;
    wire N__12245;
    wire N__12234;
    wire N__12231;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12129;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12118;
    wire N__12111;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12098;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12080;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12036;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11983;
    wire N__11978;
    wire N__11975;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11940;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11910;
    wire N__11907;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11895;
    wire N__11894;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11775;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11699;
    wire N__11694;
    wire N__11689;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11665;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11642;
    wire N__11641;
    wire N__11638;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11626;
    wire N__11623;
    wire N__11618;
    wire N__11611;
    wire N__11608;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11568;
    wire N__11567;
    wire N__11566;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11552;
    wire N__11549;
    wire N__11544;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11508;
    wire N__11505;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11493;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11477;
    wire N__11472;
    wire N__11469;
    wire N__11464;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11443;
    wire N__11440;
    wire N__11439;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11413;
    wire N__11412;
    wire N__11411;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11387;
    wire N__11380;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11358;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11352;
    wire N__11349;
    wire N__11348;
    wire N__11347;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11343;
    wire N__11340;
    wire N__11335;
    wire N__11332;
    wire N__11325;
    wire N__11316;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11205;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11189;
    wire N__11184;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11169;
    wire N__11168;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11135;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11125;
    wire N__11124;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11089;
    wire N__11084;
    wire N__11073;
    wire N__11070;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11049;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10937;
    wire N__10932;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10883;
    wire N__10878;
    wire N__10873;
    wire N__10870;
    wire N__10869;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10824;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10798;
    wire N__10795;
    wire N__10794;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10772;
    wire N__10767;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10755;
    wire N__10754;
    wire N__10751;
    wire N__10746;
    wire N__10741;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10669;
    wire N__10666;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10566;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10529;
    wire N__10524;
    wire N__10521;
    wire N__10516;
    wire N__10513;
    wire N__10512;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10488;
    wire N__10483;
    wire N__10480;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10468;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10374;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10351;
    wire N__10348;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10315;
    wire N__10306;
    wire N__10305;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10248;
    wire N__10245;
    wire N__10238;
    wire N__10235;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10206;
    wire N__10205;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10197;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10171;
    wire N__10168;
    wire N__10167;
    wire N__10166;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10146;
    wire N__10141;
    wire N__10140;
    wire N__10139;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10122;
    wire N__10117;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10103;
    wire N__10102;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10075;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10069;
    wire N__10068;
    wire N__10065;
    wire N__10056;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10011;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9945;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9923;
    wire N__9922;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9901;
    wire N__9900;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9891;
    wire N__9888;
    wire N__9883;
    wire N__9878;
    wire N__9873;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9850;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9842;
    wire N__9837;
    wire N__9832;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9813;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9799;
    wire N__9796;
    wire N__9789;
    wire N__9784;
    wire N__9783;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9731;
    wire N__9726;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9713;
    wire N__9712;
    wire N__9709;
    wire N__9702;
    wire N__9697;
    wire N__9696;
    wire N__9695;
    wire N__9692;
    wire N__9687;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9661;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9653;
    wire N__9648;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9615;
    wire N__9610;
    wire N__9607;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9589;
    wire N__9588;
    wire N__9587;
    wire N__9582;
    wire N__9579;
    wire N__9574;
    wire N__9571;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9561;
    wire N__9558;
    wire N__9553;
    wire N__9550;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9538;
    wire N__9537;
    wire N__9536;
    wire N__9535;
    wire N__9534;
    wire N__9531;
    wire N__9530;
    wire N__9521;
    wire N__9516;
    wire N__9511;
    wire N__9510;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9495;
    wire N__9494;
    wire N__9489;
    wire N__9486;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9465;
    wire N__9462;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9450;
    wire N__9445;
    wire N__9440;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9405;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9386;
    wire N__9379;
    wire N__9378;
    wire N__9377;
    wire N__9374;
    wire N__9373;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9337;
    wire N__9336;
    wire N__9333;
    wire N__9332;
    wire N__9331;
    wire N__9330;
    wire N__9327;
    wire N__9326;
    wire N__9325;
    wire N__9324;
    wire N__9323;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9317;
    wire N__9310;
    wire N__9307;
    wire N__9306;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9279;
    wire N__9276;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9212;
    wire N__9207;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9192;
    wire N__9191;
    wire N__9188;
    wire N__9183;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9171;
    wire N__9170;
    wire N__9169;
    wire N__9166;
    wire N__9161;
    wire N__9158;
    wire N__9151;
    wire N__9150;
    wire N__9149;
    wire N__9148;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9132;
    wire N__9129;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9114;
    wire N__9111;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9099;
    wire N__9098;
    wire N__9097;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9045;
    wire N__9042;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9030;
    wire N__9027;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9017;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8954;
    wire N__8949;
    wire N__8946;
    wire N__8941;
    wire N__8940;
    wire N__8939;
    wire N__8936;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8918;
    wire N__8917;
    wire N__8914;
    wire N__8909;
    wire N__8906;
    wire N__8899;
    wire N__8896;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8878;
    wire N__8877;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8863;
    wire N__8856;
    wire N__8847;
    wire N__8842;
    wire N__8835;
    wire N__8830;
    wire N__8829;
    wire N__8828;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8811;
    wire N__8806;
    wire N__8805;
    wire N__8804;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8794;
    wire N__8789;
    wire N__8782;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8760;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8742;
    wire N__8741;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8729;
    wire N__8722;
    wire N__8719;
    wire N__8718;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8668;
    wire N__8665;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8652;
    wire N__8649;
    wire N__8644;
    wire N__8643;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8631;
    wire N__8626;
    wire N__8625;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8619;
    wire N__8608;
    wire N__8605;
    wire N__8604;
    wire N__8603;
    wire N__8598;
    wire N__8595;
    wire N__8590;
    wire N__8589;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8559;
    wire N__8558;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8513;
    wire N__8508;
    wire N__8505;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8361;
    wire N__8360;
    wire N__8357;
    wire N__8356;
    wire N__8355;
    wire N__8352;
    wire N__8343;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8310;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8295;
    wire N__8294;
    wire N__8293;
    wire N__8292;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8247;
    wire N__8244;
    wire N__8237;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8211;
    wire N__8208;
    wire N__8199;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8166;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8145;
    wire N__8144;
    wire N__8143;
    wire N__8134;
    wire N__8131;
    wire N__8130;
    wire N__8127;
    wire N__8126;
    wire N__8121;
    wire N__8118;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.un143_ci_0_cascade_ ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.un4_l_count_16_cascade_ ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \buart.Z_rx.idle_0_cascade_ ;
    wire \buart.Z_rx.valid_0_cascade_ ;
    wire bu_rx_data_rdy_cascade_;
    wire \buart.Z_rx.N_27_0_i_cascade_ ;
    wire bfn_1_12_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \uu2.vbuf_count.un328_ci_3_cascade_ ;
    wire \uu2.un350_ci ;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu2.un1_l_count_2_2 ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un165_ci_0_cascade_ ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un187_ci_1 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un110_ci ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un44_ci ;
    wire \uu0.un44_ci_cascade_ ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.un66_ci ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.un88_ci_3 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un11_l_count_i ;
    wire \uu2.mem0.w_addr_0 ;
    wire \resetGen.reset_count_2_0_4 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.sample ;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_2_13_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \uu2.vbuf_raddr.un448_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.un404_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.N_34 ;
    wire \uu2.N_34_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.N_31 ;
    wire \uu2.N_31_cascade_ ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.mem0.w_data_2 ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un284_ci ;
    wire \Lab_UT.didp.countrce1.q_5_0_cascade_ ;
    wire \Lab_UT.didp.regrce3.LdAMones_0 ;
    wire G_184;
    wire G_184_cascade_;
    wire \Lab_UT.un1_idle_1_0_iclkZ0_cascade_ ;
    wire \Lab_UT.dispString.N_117_cascade_ ;
    wire G_180_cascade_;
    wire G_181_cascade_;
    wire G_180;
    wire \Lab_UT.dictrl.alarmstate_1_0_cascade_ ;
    wire G_179_cascade_;
    wire \Lab_UT.alarmstate_0_sqmuxa_1 ;
    wire \Lab_UT.un1_idle_5_0_iclkZ0_cascade_ ;
    wire \Lab_UT.un1_armed_2_0_iso_iZ0 ;
    wire G_185;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu2.un28_w_addr_user_i_cascade_ ;
    wire \uu2.un51_w_data_displaying_i_a2_1 ;
    wire \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ;
    wire \uu2.w_data_displaying_2_i_a2_i_a3_2_0 ;
    wire \INVuu2.w_addr_displaying_nesr_3C_net ;
    wire \uu2.w_addr_displaying_RNI03P31Z0Z_4 ;
    wire \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i7_mux_0 ;
    wire \uu2.N_406_cascade_ ;
    wire \uu2.bitmap_pmux ;
    wire \uu2.N_383_cascade_ ;
    wire \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ;
    wire \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ;
    wire \uu2.bitmap_pmux_u_1 ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ;
    wire \uu2.w_addr_displaying_RNI0NG56Z0Z_4 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire uart_RXD;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ;
    wire \uu2.un1_w_user_lfZ0Z_4_cascade_ ;
    wire \uu2.un20_w_addr_userZ0Z_1 ;
    wire L3_tx_data_1;
    wire L3_tx_data_4;
    wire L3_tx_data_6;
    wire \uu2.un1_w_user_lfZ0Z_3 ;
    wire \Lab_UT.dispString.N_140 ;
    wire L3_tx_data_5;
    wire G_188;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_3 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_ ;
    wire L3_tx_data_3;
    wire G_186_cascade_;
    wire G_187;
    wire G_187_cascade_;
    wire \Lab_UT.dispString.dOutP_1_iv_i_1_4 ;
    wire \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ;
    wire CONSTANT_ONE_NET;
    wire G_182;
    wire G_183;
    wire G_182_cascade_;
    wire \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ;
    wire \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.alarmstateZ0Z8 ;
    wire \Lab_UT.dictrl.g1_0_4_0_cascade_ ;
    wire \Lab_UT.dictrl.g1_0Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_5_4_0_cascade_ ;
    wire \uu2.un28_w_addr_user_i ;
    wire \INVuu2.w_addr_user_2C_net ;
    wire \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i5_mux ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.bitmap_pmux_sn_N_15_cascade_ ;
    wire \uu2.N_401 ;
    wire \INVuu2.w_addr_displaying_1_rep1_nesrC_net ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \INVuu2.bitmap_197C_net ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \Lab_UT.didp.ce_12_1 ;
    wire \Lab_UT.didp.ce_12_1_cascade_ ;
    wire \Lab_UT.didp.ce_12_3_cascade_ ;
    wire \Lab_UT.didp.countrce1.ce_12_1_1 ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_2_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_3 ;
    wire \Lab_UT.dispString.N_137 ;
    wire uu0_sec_clkD;
    wire \Lab_UT.dispString.N_143_cascade_ ;
    wire \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.dispString.un42_dOutP_1 ;
    wire \Lab_UT.dispString.N_102_cascade_ ;
    wire G_186;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_ ;
    wire L3_tx_data_2;
    wire L3_tx_data_rdy;
    wire \uu2.un1_w_user_crZ0Z_4 ;
    wire \uu2.un1_w_user_crZ0Z_3 ;
    wire G_179;
    wire G_181;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_ ;
    wire \Lab_UT.dispString.N_144 ;
    wire \Lab_UT.dispString.N_124 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_ ;
    wire \Lab_UT.dispString.N_95 ;
    wire \Lab_UT.dispString.N_102 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ;
    wire L3_tx_data_0;
    wire \Lab_UT.dispString.N_143 ;
    wire oneSecStrb;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_1 ;
    wire \Lab_UT.didp.regrce2.LdAStens_0 ;
    wire \Lab_UT.dictrl.g1_4_0 ;
    wire \Lab_UT.dictrl.g1_5_0_cascade_ ;
    wire \Lab_UT.dictrl.G_25_i_o3_3_cascade_ ;
    wire \Lab_UT.dictrl.g0_5_3_0 ;
    wire \Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ;
    wire \resetGen.escKeyZ0Z_4_cascade_ ;
    wire \resetGen.escKeyZ0 ;
    wire \resetGen.escKeyZ0Z_5 ;
    wire \Lab_UT.dictrl.g1_0Z0Z_5 ;
    wire bu_rx_data_fast_5;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ;
    wire \INVuu2.w_addr_displaying_fast_8C_net ;
    wire \uu2.N_37 ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.bitmap_pmux_sn_N_36 ;
    wire \INVuu2.bitmap_40C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \uu2.N_14_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_54_mux ;
    wire \uu2.bitmap_RNI2Q8F1Z0Z_111 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.N_24_cascade_ ;
    wire \uu2.N_31_i ;
    wire \uu2.N_166 ;
    wire \uu2.bitmap_pmux_27_ns_1_cascade_ ;
    wire \uu2.N_26 ;
    wire \uu2.N_404 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.N_149 ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.N_25 ;
    wire \Lab_UT.didp.un24_ce_3 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_ ;
    wire \Lab_UT.didp.countrce2.N_96 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_ ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_ ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ;
    wire \Lab_UT.didp.countrce4.q_5_0_cascade_ ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.didp.regrce4.LdAMtens_0 ;
    wire \Lab_UT.dispString.N_145 ;
    wire \Lab_UT.dispString.N_118_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_1 ;
    wire \Lab_UT.didp.regrce1.LdASones_0 ;
    wire \Lab_UT.dictrl.G_25_i_o3_4 ;
    wire \Lab_UT.dictrl.G_25_i_o3_5 ;
    wire \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ;
    wire \Lab_UT.dictrl.N_11_cascade_ ;
    wire \Lab_UT.dictrl.G_25_i_1_cascade_ ;
    wire \Lab_UT.dictrl.G_25_i_0 ;
    wire \Lab_UT.dictrl.G_25_i_a5_1_0 ;
    wire \Lab_UT.dictrl.N_18_0_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_6_3_0 ;
    wire \Lab_UT.dictrl.g2Z0Z_0 ;
    wire rst;
    wire \Lab_UT.dictrl.g1_1_0_0_cascade_ ;
    wire \Lab_UT.dictrl.g1_1_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1 ;
    wire \Lab_UT.dictrl.N_3 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.m37_N_2LZ0Z1 ;
    wire \Lab_UT.dictrl.N_72_mux_1 ;
    wire \Lab_UT.i8_mux_0_cascade_ ;
    wire \Lab_UT.didp.g0_0_2Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_0_sn ;
    wire \Lab_UT.dictrl.g1_1_0_1_cascade_ ;
    wire \Lab_UT.g1 ;
    wire \Lab_UT.dictrl.g0_0_rn_0 ;
    wire \Lab_UT.dictrl.m22Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_3_3_cascade_ ;
    wire \Lab_UT.dictrl.N_72_mux_0 ;
    wire bu_rx_data_fast_2;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_6;
    wire bu_rx_data_5;
    wire bu_rx_data_fast_6;
    wire \uu2.N_40 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.N_45 ;
    wire \INVuu2.w_addr_displaying_ness_6C_net ;
    wire \uu2.N_33_1 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.w_addr_7 ;
    wire o_One_Sec_Pulse;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \INVuu2.w_addr_displaying_7C_net ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.didp.reset_12_1_3 ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.startbit ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.didp.countrce2.N_93 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.un1_l_count_1_0 ;
    wire \Lab_UT.di_Stens_0 ;
    wire bu_rx_data_0;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.sec1_1 ;
    wire \Lab_UT.sec1_2 ;
    wire \Lab_UT.sec1_3 ;
    wire \Lab_UT.sec1_0 ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \uu2.bitmap_pmux_17_ns_1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.bitmap_pmux_16_ns_1 ;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_8 ;
    wire \uu2.N_44 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \Lab_UT.min2_2 ;
    wire \Lab_UT.min2_3 ;
    wire \Lab_UT.min2_0 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \INVuu2.bitmap_215C_net ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.min2_1 ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ;
    wire \Lab_UT.didp.un1_dicLdMtens_0 ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.dictrl.dicLdAMones_1 ;
    wire \Lab_UT.LdAMones ;
    wire \Lab_UT.LdAMones_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_2_fast ;
    wire \Lab_UT.dictrl.dicRun_1 ;
    wire \Lab_UT.LdASones ;
    wire \Lab_UT.LdAStens ;
    wire \Lab_UT.dictrl.N_22 ;
    wire \Lab_UT.dictrl.next_state_0_1 ;
    wire \Lab_UT.dictrl.N_20_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_22_0_0 ;
    wire \Lab_UT.didp.g0_0Z0Z_2 ;
    wire \Lab_UT.next_state_1_0_0_1_cascade_ ;
    wire \Lab_UT.dictrl.next_state6 ;
    wire \Lab_UT.dictrl.m19_1 ;
    wire \Lab_UT.dictrl.m19_1_0 ;
    wire \Lab_UT.dictrl.N_20 ;
    wire \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ;
    wire \Lab_UT.dictrl.N_20_cascade_ ;
    wire \Lab_UT.dictrl.G_14_0_a2_4_2 ;
    wire \Lab_UT.dictrl.G_14_0_0 ;
    wire \Lab_UT.dictrl.g2_0_0 ;
    wire shifter_1_rep1_RNI0FPF;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ;
    wire \Lab_UT.dictrl.G_14_0_1 ;
    wire N_15;
    wire \Lab_UT.dictrl.G_14_0_a2_1_cascade_ ;
    wire N_14_0;
    wire \Lab_UT.dictrl.N_20_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_ ;
    wire \Lab_UT.dictrl.next_state66_2 ;
    wire \Lab_UT.dictrl.state_i_3_0 ;
    wire N_5_cascade_;
    wire \Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ;
    wire \Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.N_67_mux ;
    wire \Lab_UT.dictrl.G_6_0_1_0 ;
    wire \Lab_UT.dictrl.N_12 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ;
    wire \Lab_UT.dictrl.g0_3_4 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0 ;
    wire \Lab_UT.dictrl.m22_xZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.N_72_mux_cascade_ ;
    wire bu_rx_data_4;
    wire bu_rx_data_fast_3;
    wire \Lab_UT.dictrl.m34Z0Z_1 ;
    wire \Lab_UT.dictrl.g1_0_xZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.g1_0_4 ;
    wire \Lab_UT.dictrl.g0_5_3 ;
    wire \Lab_UT.dictrl.g1_0_cascade_ ;
    wire \Lab_UT.dictrl.m22Z0Z_4 ;
    wire \Lab_UT.dictrl.g0_5Z0Z_4 ;
    wire bu_rx_data_2_rep1;
    wire bu_rx_data_0_rep1;
    wire G_6_0_a6_3_3;
    wire buart__rx_shifter_fast_4;
    wire bu_rx_data_7_rep1;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire bu_rx_data_7;
    wire \buart.Z_rx.sample_g ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.un3_w_addr_user_4_cascade_ ;
    wire \uu2.un3_w_addr_user_5 ;
    wire \uu2.un3_w_addr_user ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.un404_ci ;
    wire \uu2.un426_ci_3 ;
    wire \uu2.un404_ci_cascade_ ;
    wire \uu2.vbuf_w_addr_user.un448_ci_0 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.w_addr_user_RNI43E87Z0Z_4 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmap_pmux_20_ns_1 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.bitmap_pmux_26_bm_1 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.bitmap_RNIP2JO1Z0Z_34 ;
    wire \Lab_UT.min1_0 ;
    wire \Lab_UT.min1_3 ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmap_pmux_19_ns_1 ;
    wire \Lab_UT.sec2_0 ;
    wire \Lab_UT.sec2_3 ;
    wire \Lab_UT.sec2_1 ;
    wire \Lab_UT.sec2_2 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \uu2.bitmap_RNIM5E21Z0Z_314 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \uu2.N_152 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.didp.un1_dicLdStens_0 ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.min1_1 ;
    wire \Lab_UT.didp.countrce4.un13_qPone ;
    wire \Lab_UT.didp.countrce4.q_5_2 ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_3 ;
    wire \Lab_UT.didp.countrce1.un13_qPone_cascade_ ;
    wire \Lab_UT.loadalarm_0 ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.min1_2 ;
    wire \Lab_UT.didp.countrce1.q_5_2 ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.di_Mones_3 ;
    wire \Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.countrce4.un20_qPone ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.didp.countrce4.q_5_3 ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_1_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdMones_0 ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.state_ret_8_ess ;
    wire \Lab_UT.next_state_0 ;
    wire \Lab_UT.didp.N_90 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.LdSones_i_4 ;
    wire \Lab_UT.didp.un1_dicLdSones_0 ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.LdSones ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.didp.countrce1.q_5_1 ;
    wire \Lab_UT.dictrl.g0_1_mb_rn_0 ;
    wire \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ;
    wire \Lab_UT.dictrl.N_57_1 ;
    wire \Lab_UT.dictrl.N_55_1 ;
    wire \Lab_UT.dictrl.next_state_0_2 ;
    wire \Lab_UT.dictrl.next_state_1_2_cascade_ ;
    wire \Lab_UT.dictrl.state_i_4_2 ;
    wire \Lab_UT.bu_rx_data_rdy_0 ;
    wire \Lab_UT.dictrl.g0_1_mb_sn ;
    wire \Lab_UT.dictrl.state_i_4_1 ;
    wire \Lab_UT.dictrl.un15_loadalarm_0_cascade_ ;
    wire \Lab_UT.dictrl.loadalarm_0_0 ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire \Lab_UT.next_state_1 ;
    wire \Lab_UT.next_state_2 ;
    wire bu_rx_data_rdy;
    wire \Lab_UT.dictrl.m34_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_3 ;
    wire \Lab_UT.dictrl.next_state_1_3_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3 ;
    wire \Lab_UT.dictrl.N_33_0 ;
    wire \Lab_UT.dictrl.N_60_0_0 ;
    wire \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ;
    wire \Lab_UT.dictrl.N_26_0 ;
    wire \Lab_UT.dictrl.i8_mux_0 ;
    wire \Lab_UT.dictrl.m34_0 ;
    wire \Lab_UT.dictrl.N_18 ;
    wire \Lab_UT.dictrl.next_state_0_3 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ;
    wire \Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_ ;
    wire \Lab_UT.g0_0 ;
    wire \Lab_UT.dictrl.next_state_0_0 ;
    wire \Lab_UT.un1_next_state66_0 ;
    wire \Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ;
    wire m7_a0;
    wire \Lab_UT.dictrl.N_8_0_cascade_ ;
    wire \Lab_UT.dictrl.G_6_0_0_1_cascade_ ;
    wire \Lab_UT.dictrl.G_6_0_0 ;
    wire \Lab_UT.dictrl.N_8_0 ;
    wire \Lab_UT.dictrl.i9_mux ;
    wire \Lab_UT.dictrl.stateZ0Z_3 ;
    wire \Lab_UT.dictrl.N_60 ;
    wire \Lab_UT.dictrl.i8_mux_cascade_ ;
    wire \Lab_UT.dicLdSones_1 ;
    wire \Lab_UT.dictrl.next_state_RNO_0Z0Z_0 ;
    wire \Lab_UT.stateZ0Z_0 ;
    wire \Lab_UT.dictrl.N_59 ;
    wire bu_rx_data_3;
    wire \Lab_UT.dictrl.N_15_0 ;
    wire bu_rx_data_2;
    wire bu_rx_data_1;
    wire bu_rx_data_3_rep2;
    wire G_6_0_a6_2;
    wire \Lab_UT.dictrl.state_0_rep1 ;
    wire N_63_mux;
    wire bu_rx_data_3_rep1;
    wire \Lab_UT.dictrl.N_72_mux ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ;
    wire \Lab_UT.dictrl.m13_out ;
    wire \Lab_UT.dictrl.N_59_1_0 ;
    wire \Lab_UT.dictrl.state_fast_0 ;
    wire bu_rx_data_fast_0;
    wire bu_rx_data_fast_7;
    wire \Lab_UT.dictrl.g1_1Z0Z_5 ;
    wire bu_rx_data_1_rep1;
    wire \Lab_UT.dictrl.g1_1_4_cascade_ ;
    wire bu_rx_data_6_rep1;
    wire \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0 ;
    wire bu_rx_data_5_rep1;
    wire \Lab_UT.dictrl.g0_6_3_cascade_ ;
    wire \Lab_UT.dictrl.N_57_0 ;
    wire \Lab_UT.dictrl.g0_6_3 ;
    wire \Lab_UT.dictrl.g1_1 ;
    wire \Lab_UT.dictrl.gZ0Z2 ;
    wire Lab_UT_dictrl_state_1;
    wire \Lab_UT.dictrl.N_55_0 ;
    wire \Lab_UT.state_i_4_3 ;
    wire \Lab_UT.dictrl.g1_rn_0_cascade_ ;
    wire \Lab_UT.state_2 ;
    wire \Lab_UT.dictrl.G_25_i_a5_1_0_0 ;
    wire rst_g;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.mem0.w_addr_1 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \buart.Z_tx.un1_bitcount_c2 ;
    wire vbuf_tx_data_rdy;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.un1_bitcount_c3 ;
    wire bfn_12_2_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire clk_g;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.ser_clk ;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__8074),
            .RESETB(N__10849),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__9865,N__9850,N__9805,N__10116,N__10207,N__9832,N__9928,N__9901,N__10261}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__10417,N__13063,N__13192,N__13075,N__13123,N__16063,N__21733,N__20644,N__9247}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__9775,dangling_wire_31,N__9979,dangling_wire_32,N__9952,dangling_wire_33,N__9964,dangling_wire_34,N__10219,dangling_wire_35,N__9958,dangling_wire_36,N__9934}),
            .RCLKE(),
            .RCLK(N__22345),
            .RE(N__10845),
            .WCLKE(N__10608),
            .WCLK(N__22344),
            .WE(N__10609));
    IO_PAD led_obuft_3_iopad (
            .OE(N__22472),
            .DIN(N__22471),
            .DOUT(N__22470),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__22472),
            .PADOUT(N__22471),
            .PADIN(N__22470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__22463),
            .DIN(N__22462),
            .DOUT(N__22461),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__22463),
            .PADOUT(N__22462),
            .PADIN(N__22461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__22454),
            .DIN(N__22453),
            .DOUT(N__22452),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__22454),
            .PADOUT(N__22453),
            .PADIN(N__22452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__22445),
            .DIN(N__22444),
            .DOUT(N__22443),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__22445),
            .PADOUT(N__22444),
            .PADIN(N__22443),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__22299),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__22436),
            .DIN(N__22435),
            .DOUT(N__22434),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__22436),
            .PADOUT(N__22435),
            .PADIN(N__22434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__22427),
            .DIN(N__22426),
            .DOUT(N__22425),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__22427),
            .PADOUT(N__22426),
            .PADIN(N__22425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__22418),
            .DIN(N__22417),
            .DOUT(N__22416),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__22418),
            .PADOUT(N__22417),
            .PADIN(N__22416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__22409),
            .DIN(N__22408),
            .DOUT(N__22407),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__22409),
            .PADOUT(N__22408),
            .PADIN(N__22407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__22400),
            .DIN(N__22399),
            .DOUT(N__22398),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__22400),
            .PADOUT(N__22399),
            .PADIN(N__22398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8392),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__22391),
            .DIN(N__22390),
            .DOUT(N__22389),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__22391),
            .PADOUT(N__22390),
            .PADIN(N__22389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5450 (
            .O(N__22372),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__5449 (
            .O(N__22369),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__5448 (
            .O(N__22366),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__5447 (
            .O(N__22363),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__5446 (
            .O(N__22360),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__5445 (
            .O(N__22357),
            .I(N__22354));
    InMux I__5444 (
            .O(N__22354),
            .I(N__22351));
    LocalMux I__5443 (
            .O(N__22351),
            .I(N__22260));
    ClkMux I__5442 (
            .O(N__22350),
            .I(N__22081));
    ClkMux I__5441 (
            .O(N__22349),
            .I(N__22081));
    ClkMux I__5440 (
            .O(N__22348),
            .I(N__22081));
    ClkMux I__5439 (
            .O(N__22347),
            .I(N__22081));
    ClkMux I__5438 (
            .O(N__22346),
            .I(N__22081));
    ClkMux I__5437 (
            .O(N__22345),
            .I(N__22081));
    ClkMux I__5436 (
            .O(N__22344),
            .I(N__22081));
    ClkMux I__5435 (
            .O(N__22343),
            .I(N__22081));
    ClkMux I__5434 (
            .O(N__22342),
            .I(N__22081));
    ClkMux I__5433 (
            .O(N__22341),
            .I(N__22081));
    ClkMux I__5432 (
            .O(N__22340),
            .I(N__22081));
    ClkMux I__5431 (
            .O(N__22339),
            .I(N__22081));
    ClkMux I__5430 (
            .O(N__22338),
            .I(N__22081));
    ClkMux I__5429 (
            .O(N__22337),
            .I(N__22081));
    ClkMux I__5428 (
            .O(N__22336),
            .I(N__22081));
    ClkMux I__5427 (
            .O(N__22335),
            .I(N__22081));
    ClkMux I__5426 (
            .O(N__22334),
            .I(N__22081));
    ClkMux I__5425 (
            .O(N__22333),
            .I(N__22081));
    ClkMux I__5424 (
            .O(N__22332),
            .I(N__22081));
    ClkMux I__5423 (
            .O(N__22331),
            .I(N__22081));
    ClkMux I__5422 (
            .O(N__22330),
            .I(N__22081));
    ClkMux I__5421 (
            .O(N__22329),
            .I(N__22081));
    ClkMux I__5420 (
            .O(N__22328),
            .I(N__22081));
    ClkMux I__5419 (
            .O(N__22327),
            .I(N__22081));
    ClkMux I__5418 (
            .O(N__22326),
            .I(N__22081));
    ClkMux I__5417 (
            .O(N__22325),
            .I(N__22081));
    ClkMux I__5416 (
            .O(N__22324),
            .I(N__22081));
    ClkMux I__5415 (
            .O(N__22323),
            .I(N__22081));
    ClkMux I__5414 (
            .O(N__22322),
            .I(N__22081));
    ClkMux I__5413 (
            .O(N__22321),
            .I(N__22081));
    ClkMux I__5412 (
            .O(N__22320),
            .I(N__22081));
    ClkMux I__5411 (
            .O(N__22319),
            .I(N__22081));
    ClkMux I__5410 (
            .O(N__22318),
            .I(N__22081));
    ClkMux I__5409 (
            .O(N__22317),
            .I(N__22081));
    ClkMux I__5408 (
            .O(N__22316),
            .I(N__22081));
    ClkMux I__5407 (
            .O(N__22315),
            .I(N__22081));
    ClkMux I__5406 (
            .O(N__22314),
            .I(N__22081));
    ClkMux I__5405 (
            .O(N__22313),
            .I(N__22081));
    ClkMux I__5404 (
            .O(N__22312),
            .I(N__22081));
    ClkMux I__5403 (
            .O(N__22311),
            .I(N__22081));
    ClkMux I__5402 (
            .O(N__22310),
            .I(N__22081));
    ClkMux I__5401 (
            .O(N__22309),
            .I(N__22081));
    ClkMux I__5400 (
            .O(N__22308),
            .I(N__22081));
    ClkMux I__5399 (
            .O(N__22307),
            .I(N__22081));
    ClkMux I__5398 (
            .O(N__22306),
            .I(N__22081));
    ClkMux I__5397 (
            .O(N__22305),
            .I(N__22081));
    ClkMux I__5396 (
            .O(N__22304),
            .I(N__22081));
    ClkMux I__5395 (
            .O(N__22303),
            .I(N__22081));
    ClkMux I__5394 (
            .O(N__22302),
            .I(N__22081));
    ClkMux I__5393 (
            .O(N__22301),
            .I(N__22081));
    ClkMux I__5392 (
            .O(N__22300),
            .I(N__22081));
    ClkMux I__5391 (
            .O(N__22299),
            .I(N__22081));
    ClkMux I__5390 (
            .O(N__22298),
            .I(N__22081));
    ClkMux I__5389 (
            .O(N__22297),
            .I(N__22081));
    ClkMux I__5388 (
            .O(N__22296),
            .I(N__22081));
    ClkMux I__5387 (
            .O(N__22295),
            .I(N__22081));
    ClkMux I__5386 (
            .O(N__22294),
            .I(N__22081));
    ClkMux I__5385 (
            .O(N__22293),
            .I(N__22081));
    ClkMux I__5384 (
            .O(N__22292),
            .I(N__22081));
    ClkMux I__5383 (
            .O(N__22291),
            .I(N__22081));
    ClkMux I__5382 (
            .O(N__22290),
            .I(N__22081));
    ClkMux I__5381 (
            .O(N__22289),
            .I(N__22081));
    ClkMux I__5380 (
            .O(N__22288),
            .I(N__22081));
    ClkMux I__5379 (
            .O(N__22287),
            .I(N__22081));
    ClkMux I__5378 (
            .O(N__22286),
            .I(N__22081));
    ClkMux I__5377 (
            .O(N__22285),
            .I(N__22081));
    ClkMux I__5376 (
            .O(N__22284),
            .I(N__22081));
    ClkMux I__5375 (
            .O(N__22283),
            .I(N__22081));
    ClkMux I__5374 (
            .O(N__22282),
            .I(N__22081));
    ClkMux I__5373 (
            .O(N__22281),
            .I(N__22081));
    ClkMux I__5372 (
            .O(N__22280),
            .I(N__22081));
    ClkMux I__5371 (
            .O(N__22279),
            .I(N__22081));
    ClkMux I__5370 (
            .O(N__22278),
            .I(N__22081));
    ClkMux I__5369 (
            .O(N__22277),
            .I(N__22081));
    ClkMux I__5368 (
            .O(N__22276),
            .I(N__22081));
    ClkMux I__5367 (
            .O(N__22275),
            .I(N__22081));
    ClkMux I__5366 (
            .O(N__22274),
            .I(N__22081));
    ClkMux I__5365 (
            .O(N__22273),
            .I(N__22081));
    ClkMux I__5364 (
            .O(N__22272),
            .I(N__22081));
    ClkMux I__5363 (
            .O(N__22271),
            .I(N__22081));
    ClkMux I__5362 (
            .O(N__22270),
            .I(N__22081));
    ClkMux I__5361 (
            .O(N__22269),
            .I(N__22081));
    ClkMux I__5360 (
            .O(N__22268),
            .I(N__22081));
    ClkMux I__5359 (
            .O(N__22267),
            .I(N__22081));
    ClkMux I__5358 (
            .O(N__22266),
            .I(N__22081));
    ClkMux I__5357 (
            .O(N__22265),
            .I(N__22081));
    ClkMux I__5356 (
            .O(N__22264),
            .I(N__22081));
    ClkMux I__5355 (
            .O(N__22263),
            .I(N__22081));
    Glb2LocalMux I__5354 (
            .O(N__22260),
            .I(N__22081));
    GlobalMux I__5353 (
            .O(N__22081),
            .I(N__22078));
    gio2CtrlBuf I__5352 (
            .O(N__22078),
            .I(clk_g));
    CascadeMux I__5351 (
            .O(N__22075),
            .I(N__22072));
    InMux I__5350 (
            .O(N__22072),
            .I(N__22066));
    InMux I__5349 (
            .O(N__22071),
            .I(N__22066));
    LocalMux I__5348 (
            .O(N__22066),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__5347 (
            .O(N__22063),
            .I(N__22060));
    InMux I__5346 (
            .O(N__22060),
            .I(N__22054));
    InMux I__5345 (
            .O(N__22059),
            .I(N__22054));
    LocalMux I__5344 (
            .O(N__22054),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__5343 (
            .O(N__22051),
            .I(N__22047));
    InMux I__5342 (
            .O(N__22050),
            .I(N__22044));
    InMux I__5341 (
            .O(N__22047),
            .I(N__22041));
    LocalMux I__5340 (
            .O(N__22044),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__5339 (
            .O(N__22041),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__5338 (
            .O(N__22036),
            .I(N__22030));
    InMux I__5337 (
            .O(N__22035),
            .I(N__22030));
    LocalMux I__5336 (
            .O(N__22030),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__5335 (
            .O(N__22027),
            .I(N__22022));
    InMux I__5334 (
            .O(N__22026),
            .I(N__22017));
    InMux I__5333 (
            .O(N__22025),
            .I(N__22017));
    LocalMux I__5332 (
            .O(N__22022),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__5331 (
            .O(N__22017),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__5330 (
            .O(N__22012),
            .I(N__22007));
    InMux I__5329 (
            .O(N__22011),
            .I(N__22001));
    InMux I__5328 (
            .O(N__22010),
            .I(N__22001));
    InMux I__5327 (
            .O(N__22007),
            .I(N__21996));
    InMux I__5326 (
            .O(N__22006),
            .I(N__21996));
    LocalMux I__5325 (
            .O(N__22001),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__5324 (
            .O(N__21996),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__5323 (
            .O(N__21991),
            .I(N__21987));
    CascadeMux I__5322 (
            .O(N__21990),
            .I(N__21984));
    InMux I__5321 (
            .O(N__21987),
            .I(N__21979));
    InMux I__5320 (
            .O(N__21984),
            .I(N__21979));
    LocalMux I__5319 (
            .O(N__21979),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__5318 (
            .O(N__21976),
            .I(N__21973));
    LocalMux I__5317 (
            .O(N__21973),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    InMux I__5316 (
            .O(N__21970),
            .I(N__21960));
    InMux I__5315 (
            .O(N__21969),
            .I(N__21960));
    InMux I__5314 (
            .O(N__21968),
            .I(N__21960));
    InMux I__5313 (
            .O(N__21967),
            .I(N__21957));
    LocalMux I__5312 (
            .O(N__21960),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__5311 (
            .O(N__21957),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__5310 (
            .O(N__21952),
            .I(N__21948));
    InMux I__5309 (
            .O(N__21951),
            .I(N__21942));
    InMux I__5308 (
            .O(N__21948),
            .I(N__21935));
    InMux I__5307 (
            .O(N__21947),
            .I(N__21935));
    InMux I__5306 (
            .O(N__21946),
            .I(N__21935));
    InMux I__5305 (
            .O(N__21945),
            .I(N__21932));
    LocalMux I__5304 (
            .O(N__21942),
            .I(N__21929));
    LocalMux I__5303 (
            .O(N__21935),
            .I(N__21926));
    LocalMux I__5302 (
            .O(N__21932),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv12 I__5301 (
            .O(N__21929),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__5300 (
            .O(N__21926),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__5299 (
            .O(N__21919),
            .I(N__21914));
    InMux I__5298 (
            .O(N__21918),
            .I(N__21904));
    InMux I__5297 (
            .O(N__21917),
            .I(N__21904));
    InMux I__5296 (
            .O(N__21914),
            .I(N__21886));
    InMux I__5295 (
            .O(N__21913),
            .I(N__21886));
    InMux I__5294 (
            .O(N__21912),
            .I(N__21886));
    InMux I__5293 (
            .O(N__21911),
            .I(N__21886));
    InMux I__5292 (
            .O(N__21910),
            .I(N__21886));
    InMux I__5291 (
            .O(N__21909),
            .I(N__21886));
    LocalMux I__5290 (
            .O(N__21904),
            .I(N__21882));
    InMux I__5289 (
            .O(N__21903),
            .I(N__21879));
    InMux I__5288 (
            .O(N__21902),
            .I(N__21874));
    InMux I__5287 (
            .O(N__21901),
            .I(N__21874));
    InMux I__5286 (
            .O(N__21900),
            .I(N__21869));
    InMux I__5285 (
            .O(N__21899),
            .I(N__21869));
    LocalMux I__5284 (
            .O(N__21886),
            .I(N__21863));
    InMux I__5283 (
            .O(N__21885),
            .I(N__21860));
    Span4Mux_s2_h I__5282 (
            .O(N__21882),
            .I(N__21851));
    LocalMux I__5281 (
            .O(N__21879),
            .I(N__21851));
    LocalMux I__5280 (
            .O(N__21874),
            .I(N__21851));
    LocalMux I__5279 (
            .O(N__21869),
            .I(N__21851));
    InMux I__5278 (
            .O(N__21868),
            .I(N__21848));
    InMux I__5277 (
            .O(N__21867),
            .I(N__21845));
    InMux I__5276 (
            .O(N__21866),
            .I(N__21842));
    Span4Mux_s2_v I__5275 (
            .O(N__21863),
            .I(N__21837));
    LocalMux I__5274 (
            .O(N__21860),
            .I(N__21837));
    Span4Mux_h I__5273 (
            .O(N__21851),
            .I(N__21834));
    LocalMux I__5272 (
            .O(N__21848),
            .I(N__21831));
    LocalMux I__5271 (
            .O(N__21845),
            .I(N__21828));
    LocalMux I__5270 (
            .O(N__21842),
            .I(N__21825));
    Span4Mux_v I__5269 (
            .O(N__21837),
            .I(N__21822));
    Span4Mux_v I__5268 (
            .O(N__21834),
            .I(N__21819));
    Span4Mux_h I__5267 (
            .O(N__21831),
            .I(N__21816));
    Span4Mux_s2_v I__5266 (
            .O(N__21828),
            .I(N__21813));
    Span4Mux_s2_v I__5265 (
            .O(N__21825),
            .I(N__21810));
    Odrv4 I__5264 (
            .O(N__21822),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__5263 (
            .O(N__21819),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__5262 (
            .O(N__21816),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__5261 (
            .O(N__21813),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__5260 (
            .O(N__21810),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    InMux I__5259 (
            .O(N__21799),
            .I(N__21796));
    LocalMux I__5258 (
            .O(N__21796),
            .I(N__21793));
    Span4Mux_s1_h I__5257 (
            .O(N__21793),
            .I(N__21788));
    CascadeMux I__5256 (
            .O(N__21792),
            .I(N__21785));
    InMux I__5255 (
            .O(N__21791),
            .I(N__21777));
    Span4Mux_h I__5254 (
            .O(N__21788),
            .I(N__21770));
    InMux I__5253 (
            .O(N__21785),
            .I(N__21761));
    InMux I__5252 (
            .O(N__21784),
            .I(N__21761));
    InMux I__5251 (
            .O(N__21783),
            .I(N__21761));
    InMux I__5250 (
            .O(N__21782),
            .I(N__21761));
    InMux I__5249 (
            .O(N__21781),
            .I(N__21756));
    InMux I__5248 (
            .O(N__21780),
            .I(N__21756));
    LocalMux I__5247 (
            .O(N__21777),
            .I(N__21753));
    InMux I__5246 (
            .O(N__21776),
            .I(N__21744));
    InMux I__5245 (
            .O(N__21775),
            .I(N__21744));
    InMux I__5244 (
            .O(N__21774),
            .I(N__21744));
    InMux I__5243 (
            .O(N__21773),
            .I(N__21744));
    Odrv4 I__5242 (
            .O(N__21770),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5241 (
            .O(N__21761),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5240 (
            .O(N__21756),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__5239 (
            .O(N__21753),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5238 (
            .O(N__21744),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    CascadeMux I__5237 (
            .O(N__21733),
            .I(N__21730));
    InMux I__5236 (
            .O(N__21730),
            .I(N__21727));
    LocalMux I__5235 (
            .O(N__21727),
            .I(N__21724));
    Odrv12 I__5234 (
            .O(N__21724),
            .I(\uu2.mem0.w_addr_2 ));
    InMux I__5233 (
            .O(N__21721),
            .I(N__21718));
    LocalMux I__5232 (
            .O(N__21718),
            .I(\buart.Z_tx.un1_bitcount_c2 ));
    CascadeMux I__5231 (
            .O(N__21715),
            .I(N__21703));
    CascadeMux I__5230 (
            .O(N__21714),
            .I(N__21699));
    InMux I__5229 (
            .O(N__21713),
            .I(N__21679));
    InMux I__5228 (
            .O(N__21712),
            .I(N__21679));
    InMux I__5227 (
            .O(N__21711),
            .I(N__21679));
    InMux I__5226 (
            .O(N__21710),
            .I(N__21679));
    InMux I__5225 (
            .O(N__21709),
            .I(N__21679));
    InMux I__5224 (
            .O(N__21708),
            .I(N__21679));
    InMux I__5223 (
            .O(N__21707),
            .I(N__21679));
    InMux I__5222 (
            .O(N__21706),
            .I(N__21679));
    InMux I__5221 (
            .O(N__21703),
            .I(N__21669));
    InMux I__5220 (
            .O(N__21702),
            .I(N__21669));
    InMux I__5219 (
            .O(N__21699),
            .I(N__21669));
    InMux I__5218 (
            .O(N__21698),
            .I(N__21669));
    InMux I__5217 (
            .O(N__21697),
            .I(N__21664));
    InMux I__5216 (
            .O(N__21696),
            .I(N__21664));
    LocalMux I__5215 (
            .O(N__21679),
            .I(N__21661));
    InMux I__5214 (
            .O(N__21678),
            .I(N__21658));
    LocalMux I__5213 (
            .O(N__21669),
            .I(N__21654));
    LocalMux I__5212 (
            .O(N__21664),
            .I(N__21651));
    Span4Mux_h I__5211 (
            .O(N__21661),
            .I(N__21648));
    LocalMux I__5210 (
            .O(N__21658),
            .I(N__21645));
    InMux I__5209 (
            .O(N__21657),
            .I(N__21642));
    Span12Mux_s3_v I__5208 (
            .O(N__21654),
            .I(N__21639));
    Span4Mux_s3_v I__5207 (
            .O(N__21651),
            .I(N__21636));
    Span4Mux_h I__5206 (
            .O(N__21648),
            .I(N__21631));
    Span4Mux_s3_h I__5205 (
            .O(N__21645),
            .I(N__21631));
    LocalMux I__5204 (
            .O(N__21642),
            .I(vbuf_tx_data_rdy));
    Odrv12 I__5203 (
            .O(N__21639),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__5202 (
            .O(N__21636),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__5201 (
            .O(N__21631),
            .I(vbuf_tx_data_rdy));
    CEMux I__5200 (
            .O(N__21622),
            .I(N__21618));
    CEMux I__5199 (
            .O(N__21621),
            .I(N__21615));
    LocalMux I__5198 (
            .O(N__21618),
            .I(N__21612));
    LocalMux I__5197 (
            .O(N__21615),
            .I(N__21609));
    Span4Mux_h I__5196 (
            .O(N__21612),
            .I(N__21606));
    Span12Mux_s4_h I__5195 (
            .O(N__21609),
            .I(N__21603));
    Span4Mux_h I__5194 (
            .O(N__21606),
            .I(N__21600));
    Odrv12 I__5193 (
            .O(N__21603),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__5192 (
            .O(N__21600),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__5191 (
            .O(N__21595),
            .I(N__21591));
    InMux I__5190 (
            .O(N__21594),
            .I(N__21588));
    LocalMux I__5189 (
            .O(N__21591),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__5188 (
            .O(N__21588),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__5187 (
            .O(N__21583),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    InMux I__5186 (
            .O(N__21580),
            .I(N__21566));
    InMux I__5185 (
            .O(N__21579),
            .I(N__21566));
    InMux I__5184 (
            .O(N__21578),
            .I(N__21566));
    InMux I__5183 (
            .O(N__21577),
            .I(N__21566));
    InMux I__5182 (
            .O(N__21576),
            .I(N__21561));
    InMux I__5181 (
            .O(N__21575),
            .I(N__21561));
    LocalMux I__5180 (
            .O(N__21566),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__5179 (
            .O(N__21561),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    InMux I__5178 (
            .O(N__21556),
            .I(N__21550));
    InMux I__5177 (
            .O(N__21555),
            .I(N__21543));
    InMux I__5176 (
            .O(N__21554),
            .I(N__21543));
    InMux I__5175 (
            .O(N__21553),
            .I(N__21543));
    LocalMux I__5174 (
            .O(N__21550),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__5173 (
            .O(N__21543),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__5172 (
            .O(N__21538),
            .I(N__21535));
    InMux I__5171 (
            .O(N__21535),
            .I(N__21530));
    InMux I__5170 (
            .O(N__21534),
            .I(N__21525));
    InMux I__5169 (
            .O(N__21533),
            .I(N__21525));
    LocalMux I__5168 (
            .O(N__21530),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__5167 (
            .O(N__21525),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__5166 (
            .O(N__21520),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    InMux I__5165 (
            .O(N__21517),
            .I(N__21508));
    InMux I__5164 (
            .O(N__21516),
            .I(N__21508));
    InMux I__5163 (
            .O(N__21515),
            .I(N__21501));
    InMux I__5162 (
            .O(N__21514),
            .I(N__21501));
    InMux I__5161 (
            .O(N__21513),
            .I(N__21501));
    LocalMux I__5160 (
            .O(N__21508),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__5159 (
            .O(N__21501),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__5158 (
            .O(N__21496),
            .I(N__21493));
    LocalMux I__5157 (
            .O(N__21493),
            .I(\buart.Z_tx.un1_bitcount_c3 ));
    CascadeMux I__5156 (
            .O(N__21490),
            .I(\Lab_UT.dictrl.g0_6_3_cascade_ ));
    InMux I__5155 (
            .O(N__21487),
            .I(N__21481));
    InMux I__5154 (
            .O(N__21486),
            .I(N__21481));
    LocalMux I__5153 (
            .O(N__21481),
            .I(N__21478));
    Span4Mux_v I__5152 (
            .O(N__21478),
            .I(N__21475));
    Odrv4 I__5151 (
            .O(N__21475),
            .I(\Lab_UT.dictrl.N_57_0 ));
    InMux I__5150 (
            .O(N__21472),
            .I(N__21469));
    LocalMux I__5149 (
            .O(N__21469),
            .I(\Lab_UT.dictrl.g0_6_3 ));
    InMux I__5148 (
            .O(N__21466),
            .I(N__21460));
    InMux I__5147 (
            .O(N__21465),
            .I(N__21460));
    LocalMux I__5146 (
            .O(N__21460),
            .I(\Lab_UT.dictrl.g1_1 ));
    CascadeMux I__5145 (
            .O(N__21457),
            .I(N__21453));
    InMux I__5144 (
            .O(N__21456),
            .I(N__21448));
    InMux I__5143 (
            .O(N__21453),
            .I(N__21448));
    LocalMux I__5142 (
            .O(N__21448),
            .I(N__21445));
    Odrv12 I__5141 (
            .O(N__21445),
            .I(\Lab_UT.dictrl.gZ0Z2 ));
    InMux I__5140 (
            .O(N__21442),
            .I(N__21432));
    InMux I__5139 (
            .O(N__21441),
            .I(N__21432));
    CascadeMux I__5138 (
            .O(N__21440),
            .I(N__21420));
    InMux I__5137 (
            .O(N__21439),
            .I(N__21413));
    InMux I__5136 (
            .O(N__21438),
            .I(N__21408));
    InMux I__5135 (
            .O(N__21437),
            .I(N__21408));
    LocalMux I__5134 (
            .O(N__21432),
            .I(N__21405));
    InMux I__5133 (
            .O(N__21431),
            .I(N__21402));
    InMux I__5132 (
            .O(N__21430),
            .I(N__21393));
    InMux I__5131 (
            .O(N__21429),
            .I(N__21393));
    InMux I__5130 (
            .O(N__21428),
            .I(N__21393));
    InMux I__5129 (
            .O(N__21427),
            .I(N__21393));
    InMux I__5128 (
            .O(N__21426),
            .I(N__21390));
    InMux I__5127 (
            .O(N__21425),
            .I(N__21387));
    InMux I__5126 (
            .O(N__21424),
            .I(N__21382));
    InMux I__5125 (
            .O(N__21423),
            .I(N__21382));
    InMux I__5124 (
            .O(N__21420),
            .I(N__21377));
    InMux I__5123 (
            .O(N__21419),
            .I(N__21377));
    InMux I__5122 (
            .O(N__21418),
            .I(N__21368));
    InMux I__5121 (
            .O(N__21417),
            .I(N__21368));
    InMux I__5120 (
            .O(N__21416),
            .I(N__21365));
    LocalMux I__5119 (
            .O(N__21413),
            .I(N__21360));
    LocalMux I__5118 (
            .O(N__21408),
            .I(N__21360));
    Span4Mux_h I__5117 (
            .O(N__21405),
            .I(N__21344));
    LocalMux I__5116 (
            .O(N__21402),
            .I(N__21344));
    LocalMux I__5115 (
            .O(N__21393),
            .I(N__21344));
    LocalMux I__5114 (
            .O(N__21390),
            .I(N__21344));
    LocalMux I__5113 (
            .O(N__21387),
            .I(N__21344));
    LocalMux I__5112 (
            .O(N__21382),
            .I(N__21344));
    LocalMux I__5111 (
            .O(N__21377),
            .I(N__21344));
    InMux I__5110 (
            .O(N__21376),
            .I(N__21339));
    InMux I__5109 (
            .O(N__21375),
            .I(N__21339));
    InMux I__5108 (
            .O(N__21374),
            .I(N__21334));
    InMux I__5107 (
            .O(N__21373),
            .I(N__21334));
    LocalMux I__5106 (
            .O(N__21368),
            .I(N__21329));
    LocalMux I__5105 (
            .O(N__21365),
            .I(N__21329));
    Span4Mux_h I__5104 (
            .O(N__21360),
            .I(N__21326));
    InMux I__5103 (
            .O(N__21359),
            .I(N__21323));
    Span4Mux_v I__5102 (
            .O(N__21344),
            .I(N__21318));
    LocalMux I__5101 (
            .O(N__21339),
            .I(N__21318));
    LocalMux I__5100 (
            .O(N__21334),
            .I(Lab_UT_dictrl_state_1));
    Odrv4 I__5099 (
            .O(N__21329),
            .I(Lab_UT_dictrl_state_1));
    Odrv4 I__5098 (
            .O(N__21326),
            .I(Lab_UT_dictrl_state_1));
    LocalMux I__5097 (
            .O(N__21323),
            .I(Lab_UT_dictrl_state_1));
    Odrv4 I__5096 (
            .O(N__21318),
            .I(Lab_UT_dictrl_state_1));
    InMux I__5095 (
            .O(N__21307),
            .I(N__21304));
    LocalMux I__5094 (
            .O(N__21304),
            .I(N__21300));
    InMux I__5093 (
            .O(N__21303),
            .I(N__21297));
    Span4Mux_v I__5092 (
            .O(N__21300),
            .I(N__21294));
    LocalMux I__5091 (
            .O(N__21297),
            .I(\Lab_UT.dictrl.N_55_0 ));
    Odrv4 I__5090 (
            .O(N__21294),
            .I(\Lab_UT.dictrl.N_55_0 ));
    CascadeMux I__5089 (
            .O(N__21289),
            .I(N__21284));
    InMux I__5088 (
            .O(N__21288),
            .I(N__21279));
    InMux I__5087 (
            .O(N__21287),
            .I(N__21274));
    InMux I__5086 (
            .O(N__21284),
            .I(N__21271));
    InMux I__5085 (
            .O(N__21283),
            .I(N__21268));
    InMux I__5084 (
            .O(N__21282),
            .I(N__21265));
    LocalMux I__5083 (
            .O(N__21279),
            .I(N__21262));
    InMux I__5082 (
            .O(N__21278),
            .I(N__21259));
    CascadeMux I__5081 (
            .O(N__21277),
            .I(N__21256));
    LocalMux I__5080 (
            .O(N__21274),
            .I(N__21252));
    LocalMux I__5079 (
            .O(N__21271),
            .I(N__21247));
    LocalMux I__5078 (
            .O(N__21268),
            .I(N__21244));
    LocalMux I__5077 (
            .O(N__21265),
            .I(N__21241));
    Span4Mux_h I__5076 (
            .O(N__21262),
            .I(N__21236));
    LocalMux I__5075 (
            .O(N__21259),
            .I(N__21236));
    InMux I__5074 (
            .O(N__21256),
            .I(N__21231));
    InMux I__5073 (
            .O(N__21255),
            .I(N__21231));
    Span4Mux_h I__5072 (
            .O(N__21252),
            .I(N__21222));
    InMux I__5071 (
            .O(N__21251),
            .I(N__21219));
    InMux I__5070 (
            .O(N__21250),
            .I(N__21216));
    Span4Mux_h I__5069 (
            .O(N__21247),
            .I(N__21211));
    Span4Mux_v I__5068 (
            .O(N__21244),
            .I(N__21211));
    Span4Mux_v I__5067 (
            .O(N__21241),
            .I(N__21204));
    Span4Mux_v I__5066 (
            .O(N__21236),
            .I(N__21204));
    LocalMux I__5065 (
            .O(N__21231),
            .I(N__21204));
    InMux I__5064 (
            .O(N__21230),
            .I(N__21195));
    InMux I__5063 (
            .O(N__21229),
            .I(N__21195));
    InMux I__5062 (
            .O(N__21228),
            .I(N__21195));
    InMux I__5061 (
            .O(N__21227),
            .I(N__21195));
    InMux I__5060 (
            .O(N__21226),
            .I(N__21192));
    InMux I__5059 (
            .O(N__21225),
            .I(N__21189));
    Odrv4 I__5058 (
            .O(N__21222),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__5057 (
            .O(N__21219),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__5056 (
            .O(N__21216),
            .I(\Lab_UT.state_i_4_3 ));
    Odrv4 I__5055 (
            .O(N__21211),
            .I(\Lab_UT.state_i_4_3 ));
    Odrv4 I__5054 (
            .O(N__21204),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__5053 (
            .O(N__21195),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__5052 (
            .O(N__21192),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__5051 (
            .O(N__21189),
            .I(\Lab_UT.state_i_4_3 ));
    CascadeMux I__5050 (
            .O(N__21172),
            .I(\Lab_UT.dictrl.g1_rn_0_cascade_ ));
    InMux I__5049 (
            .O(N__21169),
            .I(N__21160));
    InMux I__5048 (
            .O(N__21168),
            .I(N__21160));
    InMux I__5047 (
            .O(N__21167),
            .I(N__21154));
    InMux I__5046 (
            .O(N__21166),
            .I(N__21154));
    InMux I__5045 (
            .O(N__21165),
            .I(N__21150));
    LocalMux I__5044 (
            .O(N__21160),
            .I(N__21147));
    InMux I__5043 (
            .O(N__21159),
            .I(N__21144));
    LocalMux I__5042 (
            .O(N__21154),
            .I(N__21136));
    InMux I__5041 (
            .O(N__21153),
            .I(N__21132));
    LocalMux I__5040 (
            .O(N__21150),
            .I(N__21129));
    Span4Mux_h I__5039 (
            .O(N__21147),
            .I(N__21126));
    LocalMux I__5038 (
            .O(N__21144),
            .I(N__21123));
    InMux I__5037 (
            .O(N__21143),
            .I(N__21120));
    InMux I__5036 (
            .O(N__21142),
            .I(N__21111));
    InMux I__5035 (
            .O(N__21141),
            .I(N__21111));
    InMux I__5034 (
            .O(N__21140),
            .I(N__21111));
    InMux I__5033 (
            .O(N__21139),
            .I(N__21111));
    Span4Mux_v I__5032 (
            .O(N__21136),
            .I(N__21103));
    InMux I__5031 (
            .O(N__21135),
            .I(N__21100));
    LocalMux I__5030 (
            .O(N__21132),
            .I(N__21097));
    Span4Mux_v I__5029 (
            .O(N__21129),
            .I(N__21092));
    Span4Mux_v I__5028 (
            .O(N__21126),
            .I(N__21092));
    Span4Mux_h I__5027 (
            .O(N__21123),
            .I(N__21085));
    LocalMux I__5026 (
            .O(N__21120),
            .I(N__21085));
    LocalMux I__5025 (
            .O(N__21111),
            .I(N__21085));
    InMux I__5024 (
            .O(N__21110),
            .I(N__21080));
    InMux I__5023 (
            .O(N__21109),
            .I(N__21080));
    InMux I__5022 (
            .O(N__21108),
            .I(N__21073));
    InMux I__5021 (
            .O(N__21107),
            .I(N__21073));
    InMux I__5020 (
            .O(N__21106),
            .I(N__21073));
    Odrv4 I__5019 (
            .O(N__21103),
            .I(\Lab_UT.state_2 ));
    LocalMux I__5018 (
            .O(N__21100),
            .I(\Lab_UT.state_2 ));
    Odrv12 I__5017 (
            .O(N__21097),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__5016 (
            .O(N__21092),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__5015 (
            .O(N__21085),
            .I(\Lab_UT.state_2 ));
    LocalMux I__5014 (
            .O(N__21080),
            .I(\Lab_UT.state_2 ));
    LocalMux I__5013 (
            .O(N__21073),
            .I(\Lab_UT.state_2 ));
    InMux I__5012 (
            .O(N__21058),
            .I(N__21055));
    LocalMux I__5011 (
            .O(N__21055),
            .I(N__21052));
    Span4Mux_h I__5010 (
            .O(N__21052),
            .I(N__21049));
    Span4Mux_v I__5009 (
            .O(N__21049),
            .I(N__21046));
    Odrv4 I__5008 (
            .O(N__21046),
            .I(\Lab_UT.dictrl.G_25_i_a5_1_0_0 ));
    CascadeMux I__5007 (
            .O(N__21043),
            .I(N__21037));
    CascadeMux I__5006 (
            .O(N__21042),
            .I(N__21029));
    CascadeMux I__5005 (
            .O(N__21041),
            .I(N__21026));
    InMux I__5004 (
            .O(N__21040),
            .I(N__21017));
    InMux I__5003 (
            .O(N__21037),
            .I(N__21014));
    InMux I__5002 (
            .O(N__21036),
            .I(N__21011));
    InMux I__5001 (
            .O(N__21035),
            .I(N__21008));
    InMux I__5000 (
            .O(N__21034),
            .I(N__21005));
    InMux I__4999 (
            .O(N__21033),
            .I(N__21002));
    InMux I__4998 (
            .O(N__21032),
            .I(N__20999));
    InMux I__4997 (
            .O(N__21029),
            .I(N__20994));
    InMux I__4996 (
            .O(N__21026),
            .I(N__20994));
    InMux I__4995 (
            .O(N__21025),
            .I(N__20989));
    InMux I__4994 (
            .O(N__21024),
            .I(N__20989));
    InMux I__4993 (
            .O(N__21023),
            .I(N__20986));
    InMux I__4992 (
            .O(N__21022),
            .I(N__20983));
    InMux I__4991 (
            .O(N__21021),
            .I(N__20978));
    InMux I__4990 (
            .O(N__21020),
            .I(N__20978));
    LocalMux I__4989 (
            .O(N__21017),
            .I(N__20975));
    LocalMux I__4988 (
            .O(N__21014),
            .I(N__20928));
    LocalMux I__4987 (
            .O(N__21011),
            .I(N__20925));
    LocalMux I__4986 (
            .O(N__21008),
            .I(N__20922));
    LocalMux I__4985 (
            .O(N__21005),
            .I(N__20919));
    LocalMux I__4984 (
            .O(N__21002),
            .I(N__20916));
    LocalMux I__4983 (
            .O(N__20999),
            .I(N__20913));
    LocalMux I__4982 (
            .O(N__20994),
            .I(N__20910));
    LocalMux I__4981 (
            .O(N__20989),
            .I(N__20907));
    LocalMux I__4980 (
            .O(N__20986),
            .I(N__20892));
    LocalMux I__4979 (
            .O(N__20983),
            .I(N__20889));
    LocalMux I__4978 (
            .O(N__20978),
            .I(N__20886));
    Glb2LocalMux I__4977 (
            .O(N__20975),
            .I(N__20749));
    SRMux I__4976 (
            .O(N__20974),
            .I(N__20749));
    SRMux I__4975 (
            .O(N__20973),
            .I(N__20749));
    SRMux I__4974 (
            .O(N__20972),
            .I(N__20749));
    SRMux I__4973 (
            .O(N__20971),
            .I(N__20749));
    SRMux I__4972 (
            .O(N__20970),
            .I(N__20749));
    SRMux I__4971 (
            .O(N__20969),
            .I(N__20749));
    SRMux I__4970 (
            .O(N__20968),
            .I(N__20749));
    SRMux I__4969 (
            .O(N__20967),
            .I(N__20749));
    SRMux I__4968 (
            .O(N__20966),
            .I(N__20749));
    SRMux I__4967 (
            .O(N__20965),
            .I(N__20749));
    SRMux I__4966 (
            .O(N__20964),
            .I(N__20749));
    SRMux I__4965 (
            .O(N__20963),
            .I(N__20749));
    SRMux I__4964 (
            .O(N__20962),
            .I(N__20749));
    SRMux I__4963 (
            .O(N__20961),
            .I(N__20749));
    SRMux I__4962 (
            .O(N__20960),
            .I(N__20749));
    SRMux I__4961 (
            .O(N__20959),
            .I(N__20749));
    SRMux I__4960 (
            .O(N__20958),
            .I(N__20749));
    SRMux I__4959 (
            .O(N__20957),
            .I(N__20749));
    SRMux I__4958 (
            .O(N__20956),
            .I(N__20749));
    SRMux I__4957 (
            .O(N__20955),
            .I(N__20749));
    SRMux I__4956 (
            .O(N__20954),
            .I(N__20749));
    SRMux I__4955 (
            .O(N__20953),
            .I(N__20749));
    SRMux I__4954 (
            .O(N__20952),
            .I(N__20749));
    SRMux I__4953 (
            .O(N__20951),
            .I(N__20749));
    SRMux I__4952 (
            .O(N__20950),
            .I(N__20749));
    SRMux I__4951 (
            .O(N__20949),
            .I(N__20749));
    SRMux I__4950 (
            .O(N__20948),
            .I(N__20749));
    SRMux I__4949 (
            .O(N__20947),
            .I(N__20749));
    SRMux I__4948 (
            .O(N__20946),
            .I(N__20749));
    SRMux I__4947 (
            .O(N__20945),
            .I(N__20749));
    SRMux I__4946 (
            .O(N__20944),
            .I(N__20749));
    SRMux I__4945 (
            .O(N__20943),
            .I(N__20749));
    SRMux I__4944 (
            .O(N__20942),
            .I(N__20749));
    SRMux I__4943 (
            .O(N__20941),
            .I(N__20749));
    SRMux I__4942 (
            .O(N__20940),
            .I(N__20749));
    SRMux I__4941 (
            .O(N__20939),
            .I(N__20749));
    SRMux I__4940 (
            .O(N__20938),
            .I(N__20749));
    SRMux I__4939 (
            .O(N__20937),
            .I(N__20749));
    SRMux I__4938 (
            .O(N__20936),
            .I(N__20749));
    SRMux I__4937 (
            .O(N__20935),
            .I(N__20749));
    SRMux I__4936 (
            .O(N__20934),
            .I(N__20749));
    SRMux I__4935 (
            .O(N__20933),
            .I(N__20749));
    SRMux I__4934 (
            .O(N__20932),
            .I(N__20749));
    SRMux I__4933 (
            .O(N__20931),
            .I(N__20749));
    Glb2LocalMux I__4932 (
            .O(N__20928),
            .I(N__20749));
    Glb2LocalMux I__4931 (
            .O(N__20925),
            .I(N__20749));
    Glb2LocalMux I__4930 (
            .O(N__20922),
            .I(N__20749));
    Glb2LocalMux I__4929 (
            .O(N__20919),
            .I(N__20749));
    Glb2LocalMux I__4928 (
            .O(N__20916),
            .I(N__20749));
    Glb2LocalMux I__4927 (
            .O(N__20913),
            .I(N__20749));
    Glb2LocalMux I__4926 (
            .O(N__20910),
            .I(N__20749));
    Glb2LocalMux I__4925 (
            .O(N__20907),
            .I(N__20749));
    SRMux I__4924 (
            .O(N__20906),
            .I(N__20749));
    SRMux I__4923 (
            .O(N__20905),
            .I(N__20749));
    SRMux I__4922 (
            .O(N__20904),
            .I(N__20749));
    SRMux I__4921 (
            .O(N__20903),
            .I(N__20749));
    SRMux I__4920 (
            .O(N__20902),
            .I(N__20749));
    SRMux I__4919 (
            .O(N__20901),
            .I(N__20749));
    SRMux I__4918 (
            .O(N__20900),
            .I(N__20749));
    SRMux I__4917 (
            .O(N__20899),
            .I(N__20749));
    SRMux I__4916 (
            .O(N__20898),
            .I(N__20749));
    SRMux I__4915 (
            .O(N__20897),
            .I(N__20749));
    SRMux I__4914 (
            .O(N__20896),
            .I(N__20749));
    SRMux I__4913 (
            .O(N__20895),
            .I(N__20749));
    Glb2LocalMux I__4912 (
            .O(N__20892),
            .I(N__20749));
    Glb2LocalMux I__4911 (
            .O(N__20889),
            .I(N__20749));
    Glb2LocalMux I__4910 (
            .O(N__20886),
            .I(N__20749));
    GlobalMux I__4909 (
            .O(N__20749),
            .I(N__20746));
    gio2CtrlBuf I__4908 (
            .O(N__20746),
            .I(rst_g));
    CascadeMux I__4907 (
            .O(N__20743),
            .I(N__20735));
    InMux I__4906 (
            .O(N__20742),
            .I(N__20732));
    InMux I__4905 (
            .O(N__20741),
            .I(N__20727));
    InMux I__4904 (
            .O(N__20740),
            .I(N__20727));
    InMux I__4903 (
            .O(N__20739),
            .I(N__20724));
    InMux I__4902 (
            .O(N__20738),
            .I(N__20719));
    InMux I__4901 (
            .O(N__20735),
            .I(N__20719));
    LocalMux I__4900 (
            .O(N__20732),
            .I(N__20716));
    LocalMux I__4899 (
            .O(N__20727),
            .I(N__20711));
    LocalMux I__4898 (
            .O(N__20724),
            .I(N__20711));
    LocalMux I__4897 (
            .O(N__20719),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv12 I__4896 (
            .O(N__20716),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__4895 (
            .O(N__20711),
            .I(\uu2.w_addr_userZ0Z_1 ));
    InMux I__4894 (
            .O(N__20704),
            .I(N__20700));
    CascadeMux I__4893 (
            .O(N__20703),
            .I(N__20697));
    LocalMux I__4892 (
            .O(N__20700),
            .I(N__20694));
    InMux I__4891 (
            .O(N__20697),
            .I(N__20691));
    Span4Mux_s1_h I__4890 (
            .O(N__20694),
            .I(N__20688));
    LocalMux I__4889 (
            .O(N__20691),
            .I(N__20674));
    Span4Mux_h I__4888 (
            .O(N__20688),
            .I(N__20674));
    InMux I__4887 (
            .O(N__20687),
            .I(N__20663));
    InMux I__4886 (
            .O(N__20686),
            .I(N__20663));
    InMux I__4885 (
            .O(N__20685),
            .I(N__20663));
    InMux I__4884 (
            .O(N__20684),
            .I(N__20663));
    InMux I__4883 (
            .O(N__20683),
            .I(N__20663));
    InMux I__4882 (
            .O(N__20682),
            .I(N__20660));
    InMux I__4881 (
            .O(N__20681),
            .I(N__20653));
    InMux I__4880 (
            .O(N__20680),
            .I(N__20653));
    InMux I__4879 (
            .O(N__20679),
            .I(N__20653));
    Odrv4 I__4878 (
            .O(N__20674),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__4877 (
            .O(N__20663),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__4876 (
            .O(N__20660),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__4875 (
            .O(N__20653),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__4874 (
            .O(N__20644),
            .I(N__20641));
    InMux I__4873 (
            .O(N__20641),
            .I(N__20638));
    LocalMux I__4872 (
            .O(N__20638),
            .I(N__20635));
    Odrv12 I__4871 (
            .O(N__20635),
            .I(\uu2.mem0.w_addr_1 ));
    InMux I__4870 (
            .O(N__20632),
            .I(N__20628));
    InMux I__4869 (
            .O(N__20631),
            .I(N__20625));
    LocalMux I__4868 (
            .O(N__20628),
            .I(N__20610));
    LocalMux I__4867 (
            .O(N__20625),
            .I(N__20607));
    InMux I__4866 (
            .O(N__20624),
            .I(N__20604));
    InMux I__4865 (
            .O(N__20623),
            .I(N__20599));
    InMux I__4864 (
            .O(N__20622),
            .I(N__20599));
    InMux I__4863 (
            .O(N__20621),
            .I(N__20596));
    InMux I__4862 (
            .O(N__20620),
            .I(N__20587));
    InMux I__4861 (
            .O(N__20619),
            .I(N__20587));
    InMux I__4860 (
            .O(N__20618),
            .I(N__20587));
    InMux I__4859 (
            .O(N__20617),
            .I(N__20587));
    InMux I__4858 (
            .O(N__20616),
            .I(N__20584));
    InMux I__4857 (
            .O(N__20615),
            .I(N__20579));
    InMux I__4856 (
            .O(N__20614),
            .I(N__20574));
    InMux I__4855 (
            .O(N__20613),
            .I(N__20574));
    Span4Mux_v I__4854 (
            .O(N__20610),
            .I(N__20569));
    Span4Mux_v I__4853 (
            .O(N__20607),
            .I(N__20569));
    LocalMux I__4852 (
            .O(N__20604),
            .I(N__20566));
    LocalMux I__4851 (
            .O(N__20599),
            .I(N__20561));
    LocalMux I__4850 (
            .O(N__20596),
            .I(N__20561));
    LocalMux I__4849 (
            .O(N__20587),
            .I(N__20556));
    LocalMux I__4848 (
            .O(N__20584),
            .I(N__20556));
    InMux I__4847 (
            .O(N__20583),
            .I(N__20553));
    InMux I__4846 (
            .O(N__20582),
            .I(N__20550));
    LocalMux I__4845 (
            .O(N__20579),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4844 (
            .O(N__20574),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4843 (
            .O(N__20569),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4842 (
            .O(N__20566),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv12 I__4841 (
            .O(N__20561),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4840 (
            .O(N__20556),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4839 (
            .O(N__20553),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4838 (
            .O(N__20550),
            .I(\Lab_UT.stateZ0Z_0 ));
    InMux I__4837 (
            .O(N__20533),
            .I(N__20527));
    InMux I__4836 (
            .O(N__20532),
            .I(N__20527));
    LocalMux I__4835 (
            .O(N__20527),
            .I(\Lab_UT.dictrl.N_59 ));
    InMux I__4834 (
            .O(N__20524),
            .I(N__20518));
    InMux I__4833 (
            .O(N__20523),
            .I(N__20512));
    InMux I__4832 (
            .O(N__20522),
            .I(N__20508));
    InMux I__4831 (
            .O(N__20521),
            .I(N__20505));
    LocalMux I__4830 (
            .O(N__20518),
            .I(N__20502));
    CascadeMux I__4829 (
            .O(N__20517),
            .I(N__20499));
    InMux I__4828 (
            .O(N__20516),
            .I(N__20495));
    InMux I__4827 (
            .O(N__20515),
            .I(N__20491));
    LocalMux I__4826 (
            .O(N__20512),
            .I(N__20488));
    InMux I__4825 (
            .O(N__20511),
            .I(N__20484));
    LocalMux I__4824 (
            .O(N__20508),
            .I(N__20478));
    LocalMux I__4823 (
            .O(N__20505),
            .I(N__20478));
    Span4Mux_v I__4822 (
            .O(N__20502),
            .I(N__20475));
    InMux I__4821 (
            .O(N__20499),
            .I(N__20470));
    InMux I__4820 (
            .O(N__20498),
            .I(N__20470));
    LocalMux I__4819 (
            .O(N__20495),
            .I(N__20465));
    InMux I__4818 (
            .O(N__20494),
            .I(N__20462));
    LocalMux I__4817 (
            .O(N__20491),
            .I(N__20456));
    Span4Mux_h I__4816 (
            .O(N__20488),
            .I(N__20453));
    InMux I__4815 (
            .O(N__20487),
            .I(N__20449));
    LocalMux I__4814 (
            .O(N__20484),
            .I(N__20446));
    CascadeMux I__4813 (
            .O(N__20483),
            .I(N__20443));
    Span4Mux_v I__4812 (
            .O(N__20478),
            .I(N__20438));
    Span4Mux_v I__4811 (
            .O(N__20475),
            .I(N__20433));
    LocalMux I__4810 (
            .O(N__20470),
            .I(N__20433));
    InMux I__4809 (
            .O(N__20469),
            .I(N__20430));
    InMux I__4808 (
            .O(N__20468),
            .I(N__20427));
    Span12Mux_s11_v I__4807 (
            .O(N__20465),
            .I(N__20422));
    LocalMux I__4806 (
            .O(N__20462),
            .I(N__20422));
    InMux I__4805 (
            .O(N__20461),
            .I(N__20419));
    InMux I__4804 (
            .O(N__20460),
            .I(N__20414));
    InMux I__4803 (
            .O(N__20459),
            .I(N__20414));
    Span4Mux_v I__4802 (
            .O(N__20456),
            .I(N__20411));
    Span4Mux_v I__4801 (
            .O(N__20453),
            .I(N__20408));
    InMux I__4800 (
            .O(N__20452),
            .I(N__20405));
    LocalMux I__4799 (
            .O(N__20449),
            .I(N__20400));
    Span4Mux_v I__4798 (
            .O(N__20446),
            .I(N__20400));
    InMux I__4797 (
            .O(N__20443),
            .I(N__20397));
    InMux I__4796 (
            .O(N__20442),
            .I(N__20392));
    InMux I__4795 (
            .O(N__20441),
            .I(N__20392));
    Span4Mux_v I__4794 (
            .O(N__20438),
            .I(N__20383));
    Span4Mux_s3_h I__4793 (
            .O(N__20433),
            .I(N__20383));
    LocalMux I__4792 (
            .O(N__20430),
            .I(N__20383));
    LocalMux I__4791 (
            .O(N__20427),
            .I(N__20383));
    Span12Mux_s4_v I__4790 (
            .O(N__20422),
            .I(N__20380));
    LocalMux I__4789 (
            .O(N__20419),
            .I(bu_rx_data_3));
    LocalMux I__4788 (
            .O(N__20414),
            .I(bu_rx_data_3));
    Odrv4 I__4787 (
            .O(N__20411),
            .I(bu_rx_data_3));
    Odrv4 I__4786 (
            .O(N__20408),
            .I(bu_rx_data_3));
    LocalMux I__4785 (
            .O(N__20405),
            .I(bu_rx_data_3));
    Odrv4 I__4784 (
            .O(N__20400),
            .I(bu_rx_data_3));
    LocalMux I__4783 (
            .O(N__20397),
            .I(bu_rx_data_3));
    LocalMux I__4782 (
            .O(N__20392),
            .I(bu_rx_data_3));
    Odrv4 I__4781 (
            .O(N__20383),
            .I(bu_rx_data_3));
    Odrv12 I__4780 (
            .O(N__20380),
            .I(bu_rx_data_3));
    InMux I__4779 (
            .O(N__20359),
            .I(N__20353));
    InMux I__4778 (
            .O(N__20358),
            .I(N__20353));
    LocalMux I__4777 (
            .O(N__20353),
            .I(N__20349));
    InMux I__4776 (
            .O(N__20352),
            .I(N__20346));
    Odrv4 I__4775 (
            .O(N__20349),
            .I(\Lab_UT.dictrl.N_15_0 ));
    LocalMux I__4774 (
            .O(N__20346),
            .I(\Lab_UT.dictrl.N_15_0 ));
    InMux I__4773 (
            .O(N__20341),
            .I(N__20331));
    InMux I__4772 (
            .O(N__20340),
            .I(N__20331));
    InMux I__4771 (
            .O(N__20339),
            .I(N__20327));
    InMux I__4770 (
            .O(N__20338),
            .I(N__20322));
    InMux I__4769 (
            .O(N__20337),
            .I(N__20319));
    InMux I__4768 (
            .O(N__20336),
            .I(N__20316));
    LocalMux I__4767 (
            .O(N__20331),
            .I(N__20313));
    InMux I__4766 (
            .O(N__20330),
            .I(N__20307));
    LocalMux I__4765 (
            .O(N__20327),
            .I(N__20304));
    InMux I__4764 (
            .O(N__20326),
            .I(N__20298));
    InMux I__4763 (
            .O(N__20325),
            .I(N__20295));
    LocalMux I__4762 (
            .O(N__20322),
            .I(N__20292));
    LocalMux I__4761 (
            .O(N__20319),
            .I(N__20287));
    LocalMux I__4760 (
            .O(N__20316),
            .I(N__20287));
    Span4Mux_v I__4759 (
            .O(N__20313),
            .I(N__20284));
    InMux I__4758 (
            .O(N__20312),
            .I(N__20279));
    InMux I__4757 (
            .O(N__20311),
            .I(N__20279));
    InMux I__4756 (
            .O(N__20310),
            .I(N__20276));
    LocalMux I__4755 (
            .O(N__20307),
            .I(N__20269));
    Sp12to4 I__4754 (
            .O(N__20304),
            .I(N__20269));
    InMux I__4753 (
            .O(N__20303),
            .I(N__20266));
    InMux I__4752 (
            .O(N__20302),
            .I(N__20263));
    CascadeMux I__4751 (
            .O(N__20301),
            .I(N__20258));
    LocalMux I__4750 (
            .O(N__20298),
            .I(N__20255));
    LocalMux I__4749 (
            .O(N__20295),
            .I(N__20248));
    Span4Mux_h I__4748 (
            .O(N__20292),
            .I(N__20248));
    Span4Mux_v I__4747 (
            .O(N__20287),
            .I(N__20248));
    Span4Mux_v I__4746 (
            .O(N__20284),
            .I(N__20241));
    LocalMux I__4745 (
            .O(N__20279),
            .I(N__20241));
    LocalMux I__4744 (
            .O(N__20276),
            .I(N__20241));
    InMux I__4743 (
            .O(N__20275),
            .I(N__20236));
    InMux I__4742 (
            .O(N__20274),
            .I(N__20236));
    Span12Mux_v I__4741 (
            .O(N__20269),
            .I(N__20233));
    LocalMux I__4740 (
            .O(N__20266),
            .I(N__20230));
    LocalMux I__4739 (
            .O(N__20263),
            .I(N__20227));
    InMux I__4738 (
            .O(N__20262),
            .I(N__20220));
    InMux I__4737 (
            .O(N__20261),
            .I(N__20220));
    InMux I__4736 (
            .O(N__20258),
            .I(N__20220));
    Span4Mux_h I__4735 (
            .O(N__20255),
            .I(N__20213));
    Span4Mux_v I__4734 (
            .O(N__20248),
            .I(N__20213));
    Span4Mux_h I__4733 (
            .O(N__20241),
            .I(N__20213));
    LocalMux I__4732 (
            .O(N__20236),
            .I(bu_rx_data_2));
    Odrv12 I__4731 (
            .O(N__20233),
            .I(bu_rx_data_2));
    Odrv4 I__4730 (
            .O(N__20230),
            .I(bu_rx_data_2));
    Odrv12 I__4729 (
            .O(N__20227),
            .I(bu_rx_data_2));
    LocalMux I__4728 (
            .O(N__20220),
            .I(bu_rx_data_2));
    Odrv4 I__4727 (
            .O(N__20213),
            .I(bu_rx_data_2));
    InMux I__4726 (
            .O(N__20200),
            .I(N__20195));
    InMux I__4725 (
            .O(N__20199),
            .I(N__20192));
    CascadeMux I__4724 (
            .O(N__20198),
            .I(N__20188));
    LocalMux I__4723 (
            .O(N__20195),
            .I(N__20178));
    LocalMux I__4722 (
            .O(N__20192),
            .I(N__20178));
    InMux I__4721 (
            .O(N__20191),
            .I(N__20174));
    InMux I__4720 (
            .O(N__20188),
            .I(N__20171));
    InMux I__4719 (
            .O(N__20187),
            .I(N__20166));
    InMux I__4718 (
            .O(N__20186),
            .I(N__20163));
    CascadeMux I__4717 (
            .O(N__20185),
            .I(N__20159));
    InMux I__4716 (
            .O(N__20184),
            .I(N__20156));
    InMux I__4715 (
            .O(N__20183),
            .I(N__20151));
    Span4Mux_v I__4714 (
            .O(N__20178),
            .I(N__20148));
    InMux I__4713 (
            .O(N__20177),
            .I(N__20145));
    LocalMux I__4712 (
            .O(N__20174),
            .I(N__20140));
    LocalMux I__4711 (
            .O(N__20171),
            .I(N__20140));
    InMux I__4710 (
            .O(N__20170),
            .I(N__20137));
    InMux I__4709 (
            .O(N__20169),
            .I(N__20134));
    LocalMux I__4708 (
            .O(N__20166),
            .I(N__20131));
    LocalMux I__4707 (
            .O(N__20163),
            .I(N__20128));
    CascadeMux I__4706 (
            .O(N__20162),
            .I(N__20123));
    InMux I__4705 (
            .O(N__20159),
            .I(N__20120));
    LocalMux I__4704 (
            .O(N__20156),
            .I(N__20117));
    InMux I__4703 (
            .O(N__20155),
            .I(N__20114));
    InMux I__4702 (
            .O(N__20154),
            .I(N__20111));
    LocalMux I__4701 (
            .O(N__20151),
            .I(N__20107));
    Span4Mux_v I__4700 (
            .O(N__20148),
            .I(N__20100));
    LocalMux I__4699 (
            .O(N__20145),
            .I(N__20100));
    Span4Mux_v I__4698 (
            .O(N__20140),
            .I(N__20100));
    LocalMux I__4697 (
            .O(N__20137),
            .I(N__20091));
    LocalMux I__4696 (
            .O(N__20134),
            .I(N__20091));
    Span4Mux_v I__4695 (
            .O(N__20131),
            .I(N__20091));
    Span4Mux_h I__4694 (
            .O(N__20128),
            .I(N__20091));
    InMux I__4693 (
            .O(N__20127),
            .I(N__20086));
    InMux I__4692 (
            .O(N__20126),
            .I(N__20086));
    InMux I__4691 (
            .O(N__20123),
            .I(N__20083));
    LocalMux I__4690 (
            .O(N__20120),
            .I(N__20080));
    Span4Mux_v I__4689 (
            .O(N__20117),
            .I(N__20077));
    LocalMux I__4688 (
            .O(N__20114),
            .I(N__20074));
    LocalMux I__4687 (
            .O(N__20111),
            .I(N__20071));
    InMux I__4686 (
            .O(N__20110),
            .I(N__20068));
    Span4Mux_h I__4685 (
            .O(N__20107),
            .I(N__20065));
    Span4Mux_h I__4684 (
            .O(N__20100),
            .I(N__20062));
    Span4Mux_v I__4683 (
            .O(N__20091),
            .I(N__20053));
    LocalMux I__4682 (
            .O(N__20086),
            .I(N__20053));
    LocalMux I__4681 (
            .O(N__20083),
            .I(N__20053));
    Span4Mux_h I__4680 (
            .O(N__20080),
            .I(N__20053));
    Odrv4 I__4679 (
            .O(N__20077),
            .I(bu_rx_data_1));
    Odrv4 I__4678 (
            .O(N__20074),
            .I(bu_rx_data_1));
    Odrv4 I__4677 (
            .O(N__20071),
            .I(bu_rx_data_1));
    LocalMux I__4676 (
            .O(N__20068),
            .I(bu_rx_data_1));
    Odrv4 I__4675 (
            .O(N__20065),
            .I(bu_rx_data_1));
    Odrv4 I__4674 (
            .O(N__20062),
            .I(bu_rx_data_1));
    Odrv4 I__4673 (
            .O(N__20053),
            .I(bu_rx_data_1));
    CascadeMux I__4672 (
            .O(N__20038),
            .I(N__20034));
    InMux I__4671 (
            .O(N__20037),
            .I(N__20025));
    InMux I__4670 (
            .O(N__20034),
            .I(N__20022));
    InMux I__4669 (
            .O(N__20033),
            .I(N__20019));
    InMux I__4668 (
            .O(N__20032),
            .I(N__20016));
    InMux I__4667 (
            .O(N__20031),
            .I(N__20011));
    InMux I__4666 (
            .O(N__20030),
            .I(N__20008));
    CascadeMux I__4665 (
            .O(N__20029),
            .I(N__20004));
    CascadeMux I__4664 (
            .O(N__20028),
            .I(N__20001));
    LocalMux I__4663 (
            .O(N__20025),
            .I(N__19998));
    LocalMux I__4662 (
            .O(N__20022),
            .I(N__19995));
    LocalMux I__4661 (
            .O(N__20019),
            .I(N__19992));
    LocalMux I__4660 (
            .O(N__20016),
            .I(N__19987));
    InMux I__4659 (
            .O(N__20015),
            .I(N__19982));
    InMux I__4658 (
            .O(N__20014),
            .I(N__19982));
    LocalMux I__4657 (
            .O(N__20011),
            .I(N__19977));
    LocalMux I__4656 (
            .O(N__20008),
            .I(N__19977));
    InMux I__4655 (
            .O(N__20007),
            .I(N__19974));
    InMux I__4654 (
            .O(N__20004),
            .I(N__19969));
    InMux I__4653 (
            .O(N__20001),
            .I(N__19969));
    Span4Mux_h I__4652 (
            .O(N__19998),
            .I(N__19966));
    Span4Mux_h I__4651 (
            .O(N__19995),
            .I(N__19961));
    Span4Mux_h I__4650 (
            .O(N__19992),
            .I(N__19961));
    InMux I__4649 (
            .O(N__19991),
            .I(N__19958));
    InMux I__4648 (
            .O(N__19990),
            .I(N__19955));
    Span4Mux_s3_v I__4647 (
            .O(N__19987),
            .I(N__19946));
    LocalMux I__4646 (
            .O(N__19982),
            .I(N__19946));
    Span4Mux_v I__4645 (
            .O(N__19977),
            .I(N__19946));
    LocalMux I__4644 (
            .O(N__19974),
            .I(N__19946));
    LocalMux I__4643 (
            .O(N__19969),
            .I(N__19943));
    Odrv4 I__4642 (
            .O(N__19966),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__4641 (
            .O(N__19961),
            .I(bu_rx_data_3_rep2));
    LocalMux I__4640 (
            .O(N__19958),
            .I(bu_rx_data_3_rep2));
    LocalMux I__4639 (
            .O(N__19955),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__4638 (
            .O(N__19946),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__4637 (
            .O(N__19943),
            .I(bu_rx_data_3_rep2));
    InMux I__4636 (
            .O(N__19930),
            .I(N__19927));
    LocalMux I__4635 (
            .O(N__19927),
            .I(N__19924));
    Odrv4 I__4634 (
            .O(N__19924),
            .I(G_6_0_a6_2));
    CascadeMux I__4633 (
            .O(N__19921),
            .I(N__19915));
    CascadeMux I__4632 (
            .O(N__19920),
            .I(N__19912));
    CascadeMux I__4631 (
            .O(N__19919),
            .I(N__19909));
    InMux I__4630 (
            .O(N__19918),
            .I(N__19902));
    InMux I__4629 (
            .O(N__19915),
            .I(N__19899));
    InMux I__4628 (
            .O(N__19912),
            .I(N__19896));
    InMux I__4627 (
            .O(N__19909),
            .I(N__19891));
    InMux I__4626 (
            .O(N__19908),
            .I(N__19886));
    InMux I__4625 (
            .O(N__19907),
            .I(N__19886));
    InMux I__4624 (
            .O(N__19906),
            .I(N__19881));
    InMux I__4623 (
            .O(N__19905),
            .I(N__19881));
    LocalMux I__4622 (
            .O(N__19902),
            .I(N__19876));
    LocalMux I__4621 (
            .O(N__19899),
            .I(N__19876));
    LocalMux I__4620 (
            .O(N__19896),
            .I(N__19873));
    InMux I__4619 (
            .O(N__19895),
            .I(N__19870));
    InMux I__4618 (
            .O(N__19894),
            .I(N__19865));
    LocalMux I__4617 (
            .O(N__19891),
            .I(N__19852));
    LocalMux I__4616 (
            .O(N__19886),
            .I(N__19852));
    LocalMux I__4615 (
            .O(N__19881),
            .I(N__19852));
    Span4Mux_h I__4614 (
            .O(N__19876),
            .I(N__19852));
    Span4Mux_h I__4613 (
            .O(N__19873),
            .I(N__19852));
    LocalMux I__4612 (
            .O(N__19870),
            .I(N__19852));
    InMux I__4611 (
            .O(N__19869),
            .I(N__19849));
    InMux I__4610 (
            .O(N__19868),
            .I(N__19846));
    LocalMux I__4609 (
            .O(N__19865),
            .I(N__19843));
    Span4Mux_v I__4608 (
            .O(N__19852),
            .I(N__19840));
    LocalMux I__4607 (
            .O(N__19849),
            .I(N__19835));
    LocalMux I__4606 (
            .O(N__19846),
            .I(N__19835));
    Odrv4 I__4605 (
            .O(N__19843),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv4 I__4604 (
            .O(N__19840),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv12 I__4603 (
            .O(N__19835),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    InMux I__4602 (
            .O(N__19828),
            .I(N__19811));
    InMux I__4601 (
            .O(N__19827),
            .I(N__19811));
    InMux I__4600 (
            .O(N__19826),
            .I(N__19808));
    InMux I__4599 (
            .O(N__19825),
            .I(N__19801));
    InMux I__4598 (
            .O(N__19824),
            .I(N__19801));
    InMux I__4597 (
            .O(N__19823),
            .I(N__19801));
    InMux I__4596 (
            .O(N__19822),
            .I(N__19795));
    InMux I__4595 (
            .O(N__19821),
            .I(N__19795));
    InMux I__4594 (
            .O(N__19820),
            .I(N__19790));
    InMux I__4593 (
            .O(N__19819),
            .I(N__19790));
    InMux I__4592 (
            .O(N__19818),
            .I(N__19783));
    InMux I__4591 (
            .O(N__19817),
            .I(N__19783));
    InMux I__4590 (
            .O(N__19816),
            .I(N__19783));
    LocalMux I__4589 (
            .O(N__19811),
            .I(N__19780));
    LocalMux I__4588 (
            .O(N__19808),
            .I(N__19773));
    LocalMux I__4587 (
            .O(N__19801),
            .I(N__19773));
    InMux I__4586 (
            .O(N__19800),
            .I(N__19770));
    LocalMux I__4585 (
            .O(N__19795),
            .I(N__19767));
    LocalMux I__4584 (
            .O(N__19790),
            .I(N__19762));
    LocalMux I__4583 (
            .O(N__19783),
            .I(N__19762));
    Span4Mux_h I__4582 (
            .O(N__19780),
            .I(N__19759));
    InMux I__4581 (
            .O(N__19779),
            .I(N__19754));
    InMux I__4580 (
            .O(N__19778),
            .I(N__19754));
    Span4Mux_v I__4579 (
            .O(N__19773),
            .I(N__19751));
    LocalMux I__4578 (
            .O(N__19770),
            .I(N_63_mux));
    Odrv4 I__4577 (
            .O(N__19767),
            .I(N_63_mux));
    Odrv4 I__4576 (
            .O(N__19762),
            .I(N_63_mux));
    Odrv4 I__4575 (
            .O(N__19759),
            .I(N_63_mux));
    LocalMux I__4574 (
            .O(N__19754),
            .I(N_63_mux));
    Odrv4 I__4573 (
            .O(N__19751),
            .I(N_63_mux));
    CascadeMux I__4572 (
            .O(N__19738),
            .I(N__19732));
    CascadeMux I__4571 (
            .O(N__19737),
            .I(N__19727));
    CascadeMux I__4570 (
            .O(N__19736),
            .I(N__19724));
    InMux I__4569 (
            .O(N__19735),
            .I(N__19720));
    InMux I__4568 (
            .O(N__19732),
            .I(N__19715));
    InMux I__4567 (
            .O(N__19731),
            .I(N__19715));
    CascadeMux I__4566 (
            .O(N__19730),
            .I(N__19710));
    InMux I__4565 (
            .O(N__19727),
            .I(N__19707));
    InMux I__4564 (
            .O(N__19724),
            .I(N__19704));
    CascadeMux I__4563 (
            .O(N__19723),
            .I(N__19701));
    LocalMux I__4562 (
            .O(N__19720),
            .I(N__19696));
    LocalMux I__4561 (
            .O(N__19715),
            .I(N__19696));
    InMux I__4560 (
            .O(N__19714),
            .I(N__19692));
    InMux I__4559 (
            .O(N__19713),
            .I(N__19688));
    InMux I__4558 (
            .O(N__19710),
            .I(N__19685));
    LocalMux I__4557 (
            .O(N__19707),
            .I(N__19680));
    LocalMux I__4556 (
            .O(N__19704),
            .I(N__19680));
    InMux I__4555 (
            .O(N__19701),
            .I(N__19677));
    Span4Mux_v I__4554 (
            .O(N__19696),
            .I(N__19674));
    InMux I__4553 (
            .O(N__19695),
            .I(N__19671));
    LocalMux I__4552 (
            .O(N__19692),
            .I(N__19668));
    InMux I__4551 (
            .O(N__19691),
            .I(N__19665));
    LocalMux I__4550 (
            .O(N__19688),
            .I(N__19656));
    LocalMux I__4549 (
            .O(N__19685),
            .I(N__19656));
    Span4Mux_v I__4548 (
            .O(N__19680),
            .I(N__19656));
    LocalMux I__4547 (
            .O(N__19677),
            .I(N__19656));
    Span4Mux_s2_v I__4546 (
            .O(N__19674),
            .I(N__19653));
    LocalMux I__4545 (
            .O(N__19671),
            .I(N__19646));
    Span4Mux_v I__4544 (
            .O(N__19668),
            .I(N__19646));
    LocalMux I__4543 (
            .O(N__19665),
            .I(N__19646));
    Span4Mux_h I__4542 (
            .O(N__19656),
            .I(N__19643));
    Odrv4 I__4541 (
            .O(N__19653),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__4540 (
            .O(N__19646),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__4539 (
            .O(N__19643),
            .I(bu_rx_data_3_rep1));
    InMux I__4538 (
            .O(N__19636),
            .I(N__19633));
    LocalMux I__4537 (
            .O(N__19633),
            .I(N__19628));
    InMux I__4536 (
            .O(N__19632),
            .I(N__19624));
    InMux I__4535 (
            .O(N__19631),
            .I(N__19621));
    Span4Mux_h I__4534 (
            .O(N__19628),
            .I(N__19618));
    InMux I__4533 (
            .O(N__19627),
            .I(N__19615));
    LocalMux I__4532 (
            .O(N__19624),
            .I(\Lab_UT.dictrl.N_72_mux ));
    LocalMux I__4531 (
            .O(N__19621),
            .I(\Lab_UT.dictrl.N_72_mux ));
    Odrv4 I__4530 (
            .O(N__19618),
            .I(\Lab_UT.dictrl.N_72_mux ));
    LocalMux I__4529 (
            .O(N__19615),
            .I(\Lab_UT.dictrl.N_72_mux ));
    InMux I__4528 (
            .O(N__19606),
            .I(N__19603));
    LocalMux I__4527 (
            .O(N__19603),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ));
    CascadeMux I__4526 (
            .O(N__19600),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ));
    InMux I__4525 (
            .O(N__19597),
            .I(N__19591));
    InMux I__4524 (
            .O(N__19596),
            .I(N__19591));
    LocalMux I__4523 (
            .O(N__19591),
            .I(N__19584));
    InMux I__4522 (
            .O(N__19590),
            .I(N__19579));
    InMux I__4521 (
            .O(N__19589),
            .I(N__19579));
    InMux I__4520 (
            .O(N__19588),
            .I(N__19575));
    InMux I__4519 (
            .O(N__19587),
            .I(N__19572));
    Span4Mux_v I__4518 (
            .O(N__19584),
            .I(N__19567));
    LocalMux I__4517 (
            .O(N__19579),
            .I(N__19567));
    InMux I__4516 (
            .O(N__19578),
            .I(N__19564));
    LocalMux I__4515 (
            .O(N__19575),
            .I(\Lab_UT.dictrl.m13_out ));
    LocalMux I__4514 (
            .O(N__19572),
            .I(\Lab_UT.dictrl.m13_out ));
    Odrv4 I__4513 (
            .O(N__19567),
            .I(\Lab_UT.dictrl.m13_out ));
    LocalMux I__4512 (
            .O(N__19564),
            .I(\Lab_UT.dictrl.m13_out ));
    InMux I__4511 (
            .O(N__19555),
            .I(N__19552));
    LocalMux I__4510 (
            .O(N__19552),
            .I(N__19549));
    Odrv12 I__4509 (
            .O(N__19549),
            .I(\Lab_UT.dictrl.N_59_1_0 ));
    InMux I__4508 (
            .O(N__19546),
            .I(N__19541));
    CascadeMux I__4507 (
            .O(N__19545),
            .I(N__19538));
    CascadeMux I__4506 (
            .O(N__19544),
            .I(N__19535));
    LocalMux I__4505 (
            .O(N__19541),
            .I(N__19532));
    InMux I__4504 (
            .O(N__19538),
            .I(N__19529));
    InMux I__4503 (
            .O(N__19535),
            .I(N__19526));
    Span4Mux_v I__4502 (
            .O(N__19532),
            .I(N__19523));
    LocalMux I__4501 (
            .O(N__19529),
            .I(N__19518));
    LocalMux I__4500 (
            .O(N__19526),
            .I(N__19518));
    Odrv4 I__4499 (
            .O(N__19523),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    Odrv12 I__4498 (
            .O(N__19518),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    InMux I__4497 (
            .O(N__19513),
            .I(N__19509));
    InMux I__4496 (
            .O(N__19512),
            .I(N__19506));
    LocalMux I__4495 (
            .O(N__19509),
            .I(N__19503));
    LocalMux I__4494 (
            .O(N__19506),
            .I(bu_rx_data_fast_0));
    Odrv4 I__4493 (
            .O(N__19503),
            .I(bu_rx_data_fast_0));
    InMux I__4492 (
            .O(N__19498),
            .I(N__19495));
    LocalMux I__4491 (
            .O(N__19495),
            .I(N__19491));
    CascadeMux I__4490 (
            .O(N__19494),
            .I(N__19488));
    Span4Mux_h I__4489 (
            .O(N__19491),
            .I(N__19485));
    InMux I__4488 (
            .O(N__19488),
            .I(N__19482));
    Odrv4 I__4487 (
            .O(N__19485),
            .I(bu_rx_data_fast_7));
    LocalMux I__4486 (
            .O(N__19482),
            .I(bu_rx_data_fast_7));
    InMux I__4485 (
            .O(N__19477),
            .I(N__19474));
    LocalMux I__4484 (
            .O(N__19474),
            .I(N__19471));
    Span4Mux_s3_h I__4483 (
            .O(N__19471),
            .I(N__19468));
    Odrv4 I__4482 (
            .O(N__19468),
            .I(\Lab_UT.dictrl.g1_1Z0Z_5 ));
    InMux I__4481 (
            .O(N__19465),
            .I(N__19461));
    InMux I__4480 (
            .O(N__19464),
            .I(N__19458));
    LocalMux I__4479 (
            .O(N__19461),
            .I(N__19446));
    LocalMux I__4478 (
            .O(N__19458),
            .I(N__19446));
    InMux I__4477 (
            .O(N__19457),
            .I(N__19443));
    InMux I__4476 (
            .O(N__19456),
            .I(N__19438));
    InMux I__4475 (
            .O(N__19455),
            .I(N__19438));
    InMux I__4474 (
            .O(N__19454),
            .I(N__19435));
    InMux I__4473 (
            .O(N__19453),
            .I(N__19430));
    InMux I__4472 (
            .O(N__19452),
            .I(N__19430));
    InMux I__4471 (
            .O(N__19451),
            .I(N__19427));
    Span4Mux_h I__4470 (
            .O(N__19446),
            .I(N__19420));
    LocalMux I__4469 (
            .O(N__19443),
            .I(N__19420));
    LocalMux I__4468 (
            .O(N__19438),
            .I(N__19420));
    LocalMux I__4467 (
            .O(N__19435),
            .I(N__19417));
    LocalMux I__4466 (
            .O(N__19430),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4465 (
            .O(N__19427),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__4464 (
            .O(N__19420),
            .I(bu_rx_data_1_rep1));
    Odrv12 I__4463 (
            .O(N__19417),
            .I(bu_rx_data_1_rep1));
    CascadeMux I__4462 (
            .O(N__19408),
            .I(\Lab_UT.dictrl.g1_1_4_cascade_ ));
    CascadeMux I__4461 (
            .O(N__19405),
            .I(N__19400));
    InMux I__4460 (
            .O(N__19404),
            .I(N__19395));
    InMux I__4459 (
            .O(N__19403),
            .I(N__19392));
    InMux I__4458 (
            .O(N__19400),
            .I(N__19385));
    InMux I__4457 (
            .O(N__19399),
            .I(N__19385));
    InMux I__4456 (
            .O(N__19398),
            .I(N__19385));
    LocalMux I__4455 (
            .O(N__19395),
            .I(bu_rx_data_6_rep1));
    LocalMux I__4454 (
            .O(N__19392),
            .I(bu_rx_data_6_rep1));
    LocalMux I__4453 (
            .O(N__19385),
            .I(bu_rx_data_6_rep1));
    InMux I__4452 (
            .O(N__19378),
            .I(N__19375));
    LocalMux I__4451 (
            .O(N__19375),
            .I(\Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0 ));
    InMux I__4450 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__4449 (
            .O(N__19369),
            .I(N__19366));
    Span4Mux_v I__4448 (
            .O(N__19366),
            .I(N__19360));
    InMux I__4447 (
            .O(N__19365),
            .I(N__19357));
    InMux I__4446 (
            .O(N__19364),
            .I(N__19352));
    InMux I__4445 (
            .O(N__19363),
            .I(N__19352));
    Odrv4 I__4444 (
            .O(N__19360),
            .I(bu_rx_data_5_rep1));
    LocalMux I__4443 (
            .O(N__19357),
            .I(bu_rx_data_5_rep1));
    LocalMux I__4442 (
            .O(N__19352),
            .I(bu_rx_data_5_rep1));
    CascadeMux I__4441 (
            .O(N__19345),
            .I(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_ ));
    CEMux I__4440 (
            .O(N__19342),
            .I(N__19338));
    CEMux I__4439 (
            .O(N__19341),
            .I(N__19335));
    LocalMux I__4438 (
            .O(N__19338),
            .I(N__19332));
    LocalMux I__4437 (
            .O(N__19335),
            .I(N__19328));
    Span4Mux_v I__4436 (
            .O(N__19332),
            .I(N__19324));
    CEMux I__4435 (
            .O(N__19331),
            .I(N__19321));
    Span4Mux_v I__4434 (
            .O(N__19328),
            .I(N__19318));
    CEMux I__4433 (
            .O(N__19327),
            .I(N__19315));
    Span4Mux_v I__4432 (
            .O(N__19324),
            .I(N__19310));
    LocalMux I__4431 (
            .O(N__19321),
            .I(N__19310));
    Span4Mux_s2_h I__4430 (
            .O(N__19318),
            .I(N__19307));
    LocalMux I__4429 (
            .O(N__19315),
            .I(N__19304));
    Span4Mux_h I__4428 (
            .O(N__19310),
            .I(N__19301));
    Odrv4 I__4427 (
            .O(N__19307),
            .I(\Lab_UT.g0_0 ));
    Odrv12 I__4426 (
            .O(N__19304),
            .I(\Lab_UT.g0_0 ));
    Odrv4 I__4425 (
            .O(N__19301),
            .I(\Lab_UT.g0_0 ));
    CascadeMux I__4424 (
            .O(N__19294),
            .I(N__19291));
    InMux I__4423 (
            .O(N__19291),
            .I(N__19287));
    InMux I__4422 (
            .O(N__19290),
            .I(N__19284));
    LocalMux I__4421 (
            .O(N__19287),
            .I(N__19281));
    LocalMux I__4420 (
            .O(N__19284),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    Odrv4 I__4419 (
            .O(N__19281),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    CascadeMux I__4418 (
            .O(N__19276),
            .I(N__19271));
    CascadeMux I__4417 (
            .O(N__19275),
            .I(N__19268));
    CascadeMux I__4416 (
            .O(N__19274),
            .I(N__19260));
    InMux I__4415 (
            .O(N__19271),
            .I(N__19247));
    InMux I__4414 (
            .O(N__19268),
            .I(N__19247));
    InMux I__4413 (
            .O(N__19267),
            .I(N__19247));
    InMux I__4412 (
            .O(N__19266),
            .I(N__19247));
    InMux I__4411 (
            .O(N__19265),
            .I(N__19239));
    InMux I__4410 (
            .O(N__19264),
            .I(N__19239));
    InMux I__4409 (
            .O(N__19263),
            .I(N__19232));
    InMux I__4408 (
            .O(N__19260),
            .I(N__19232));
    InMux I__4407 (
            .O(N__19259),
            .I(N__19232));
    InMux I__4406 (
            .O(N__19258),
            .I(N__19219));
    InMux I__4405 (
            .O(N__19257),
            .I(N__19219));
    InMux I__4404 (
            .O(N__19256),
            .I(N__19219));
    LocalMux I__4403 (
            .O(N__19247),
            .I(N__19216));
    InMux I__4402 (
            .O(N__19246),
            .I(N__19213));
    CascadeMux I__4401 (
            .O(N__19245),
            .I(N__19210));
    InMux I__4400 (
            .O(N__19244),
            .I(N__19205));
    LocalMux I__4399 (
            .O(N__19239),
            .I(N__19202));
    LocalMux I__4398 (
            .O(N__19232),
            .I(N__19199));
    InMux I__4397 (
            .O(N__19231),
            .I(N__19192));
    InMux I__4396 (
            .O(N__19230),
            .I(N__19192));
    InMux I__4395 (
            .O(N__19229),
            .I(N__19192));
    InMux I__4394 (
            .O(N__19228),
            .I(N__19187));
    InMux I__4393 (
            .O(N__19227),
            .I(N__19187));
    InMux I__4392 (
            .O(N__19226),
            .I(N__19184));
    LocalMux I__4391 (
            .O(N__19219),
            .I(N__19181));
    Span4Mux_v I__4390 (
            .O(N__19216),
            .I(N__19176));
    LocalMux I__4389 (
            .O(N__19213),
            .I(N__19176));
    InMux I__4388 (
            .O(N__19210),
            .I(N__19173));
    InMux I__4387 (
            .O(N__19209),
            .I(N__19168));
    InMux I__4386 (
            .O(N__19208),
            .I(N__19168));
    LocalMux I__4385 (
            .O(N__19205),
            .I(N__19161));
    Span4Mux_v I__4384 (
            .O(N__19202),
            .I(N__19161));
    Span4Mux_v I__4383 (
            .O(N__19199),
            .I(N__19161));
    LocalMux I__4382 (
            .O(N__19192),
            .I(N__19158));
    LocalMux I__4381 (
            .O(N__19187),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4380 (
            .O(N__19184),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv4 I__4379 (
            .O(N__19181),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv4 I__4378 (
            .O(N__19176),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4377 (
            .O(N__19173),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4376 (
            .O(N__19168),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv4 I__4375 (
            .O(N__19161),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv12 I__4374 (
            .O(N__19158),
            .I(\Lab_UT.un1_next_state66_0 ));
    CascadeMux I__4373 (
            .O(N__19141),
            .I(\Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ));
    InMux I__4372 (
            .O(N__19138),
            .I(N__19132));
    InMux I__4371 (
            .O(N__19137),
            .I(N__19132));
    LocalMux I__4370 (
            .O(N__19132),
            .I(N__19129));
    Span4Mux_h I__4369 (
            .O(N__19129),
            .I(N__19126));
    Odrv4 I__4368 (
            .O(N__19126),
            .I(\Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ));
    InMux I__4367 (
            .O(N__19123),
            .I(N__19118));
    InMux I__4366 (
            .O(N__19122),
            .I(N__19113));
    InMux I__4365 (
            .O(N__19121),
            .I(N__19113));
    LocalMux I__4364 (
            .O(N__19118),
            .I(N__19107));
    LocalMux I__4363 (
            .O(N__19113),
            .I(N__19107));
    InMux I__4362 (
            .O(N__19112),
            .I(N__19104));
    Span4Mux_h I__4361 (
            .O(N__19107),
            .I(N__19101));
    LocalMux I__4360 (
            .O(N__19104),
            .I(m7_a0));
    Odrv4 I__4359 (
            .O(N__19101),
            .I(m7_a0));
    CascadeMux I__4358 (
            .O(N__19096),
            .I(\Lab_UT.dictrl.N_8_0_cascade_ ));
    CascadeMux I__4357 (
            .O(N__19093),
            .I(\Lab_UT.dictrl.G_6_0_0_1_cascade_ ));
    InMux I__4356 (
            .O(N__19090),
            .I(N__19087));
    LocalMux I__4355 (
            .O(N__19087),
            .I(\Lab_UT.dictrl.G_6_0_0 ));
    InMux I__4354 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__4353 (
            .O(N__19081),
            .I(\Lab_UT.dictrl.N_8_0 ));
    InMux I__4352 (
            .O(N__19078),
            .I(N__19075));
    LocalMux I__4351 (
            .O(N__19075),
            .I(\Lab_UT.dictrl.i9_mux ));
    CascadeMux I__4350 (
            .O(N__19072),
            .I(N__19065));
    CascadeMux I__4349 (
            .O(N__19071),
            .I(N__19058));
    InMux I__4348 (
            .O(N__19070),
            .I(N__19055));
    InMux I__4347 (
            .O(N__19069),
            .I(N__19042));
    InMux I__4346 (
            .O(N__19068),
            .I(N__19042));
    InMux I__4345 (
            .O(N__19065),
            .I(N__19042));
    InMux I__4344 (
            .O(N__19064),
            .I(N__19035));
    InMux I__4343 (
            .O(N__19063),
            .I(N__19035));
    InMux I__4342 (
            .O(N__19062),
            .I(N__19035));
    InMux I__4341 (
            .O(N__19061),
            .I(N__19031));
    InMux I__4340 (
            .O(N__19058),
            .I(N__19027));
    LocalMux I__4339 (
            .O(N__19055),
            .I(N__19024));
    InMux I__4338 (
            .O(N__19054),
            .I(N__19021));
    InMux I__4337 (
            .O(N__19053),
            .I(N__19018));
    InMux I__4336 (
            .O(N__19052),
            .I(N__19015));
    InMux I__4335 (
            .O(N__19051),
            .I(N__19008));
    InMux I__4334 (
            .O(N__19050),
            .I(N__19008));
    InMux I__4333 (
            .O(N__19049),
            .I(N__19008));
    LocalMux I__4332 (
            .O(N__19042),
            .I(N__19003));
    LocalMux I__4331 (
            .O(N__19035),
            .I(N__19003));
    InMux I__4330 (
            .O(N__19034),
            .I(N__19000));
    LocalMux I__4329 (
            .O(N__19031),
            .I(N__18997));
    InMux I__4328 (
            .O(N__19030),
            .I(N__18994));
    LocalMux I__4327 (
            .O(N__19027),
            .I(N__18989));
    Span4Mux_v I__4326 (
            .O(N__19024),
            .I(N__18989));
    LocalMux I__4325 (
            .O(N__19021),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4324 (
            .O(N__19018),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4323 (
            .O(N__19015),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4322 (
            .O(N__19008),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4321 (
            .O(N__19003),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4320 (
            .O(N__19000),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4319 (
            .O(N__18997),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4318 (
            .O(N__18994),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4317 (
            .O(N__18989),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    CascadeMux I__4316 (
            .O(N__18970),
            .I(N__18966));
    InMux I__4315 (
            .O(N__18969),
            .I(N__18962));
    InMux I__4314 (
            .O(N__18966),
            .I(N__18957));
    InMux I__4313 (
            .O(N__18965),
            .I(N__18957));
    LocalMux I__4312 (
            .O(N__18962),
            .I(\Lab_UT.dictrl.N_60 ));
    LocalMux I__4311 (
            .O(N__18957),
            .I(\Lab_UT.dictrl.N_60 ));
    CascadeMux I__4310 (
            .O(N__18952),
            .I(\Lab_UT.dictrl.i8_mux_cascade_ ));
    CascadeMux I__4309 (
            .O(N__18949),
            .I(N__18945));
    InMux I__4308 (
            .O(N__18948),
            .I(N__18942));
    InMux I__4307 (
            .O(N__18945),
            .I(N__18939));
    LocalMux I__4306 (
            .O(N__18942),
            .I(N__18932));
    LocalMux I__4305 (
            .O(N__18939),
            .I(N__18929));
    InMux I__4304 (
            .O(N__18938),
            .I(N__18924));
    InMux I__4303 (
            .O(N__18937),
            .I(N__18924));
    InMux I__4302 (
            .O(N__18936),
            .I(N__18921));
    InMux I__4301 (
            .O(N__18935),
            .I(N__18917));
    Span4Mux_v I__4300 (
            .O(N__18932),
            .I(N__18914));
    Span4Mux_h I__4299 (
            .O(N__18929),
            .I(N__18907));
    LocalMux I__4298 (
            .O(N__18924),
            .I(N__18907));
    LocalMux I__4297 (
            .O(N__18921),
            .I(N__18907));
    InMux I__4296 (
            .O(N__18920),
            .I(N__18904));
    LocalMux I__4295 (
            .O(N__18917),
            .I(\Lab_UT.dicLdSones_1 ));
    Odrv4 I__4294 (
            .O(N__18914),
            .I(\Lab_UT.dicLdSones_1 ));
    Odrv4 I__4293 (
            .O(N__18907),
            .I(\Lab_UT.dicLdSones_1 ));
    LocalMux I__4292 (
            .O(N__18904),
            .I(\Lab_UT.dicLdSones_1 ));
    InMux I__4291 (
            .O(N__18895),
            .I(N__18892));
    LocalMux I__4290 (
            .O(N__18892),
            .I(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0 ));
    CascadeMux I__4289 (
            .O(N__18889),
            .I(\Lab_UT.dictrl.m34_0_cascade_ ));
    InMux I__4288 (
            .O(N__18886),
            .I(N__18883));
    LocalMux I__4287 (
            .O(N__18883),
            .I(N__18880));
    Span4Mux_v I__4286 (
            .O(N__18880),
            .I(N__18875));
    InMux I__4285 (
            .O(N__18879),
            .I(N__18870));
    InMux I__4284 (
            .O(N__18878),
            .I(N__18870));
    Odrv4 I__4283 (
            .O(N__18875),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    LocalMux I__4282 (
            .O(N__18870),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    CascadeMux I__4281 (
            .O(N__18865),
            .I(\Lab_UT.dictrl.next_state_1_3_cascade_ ));
    CascadeMux I__4280 (
            .O(N__18862),
            .I(N__18858));
    CascadeMux I__4279 (
            .O(N__18861),
            .I(N__18854));
    InMux I__4278 (
            .O(N__18858),
            .I(N__18847));
    InMux I__4277 (
            .O(N__18857),
            .I(N__18847));
    InMux I__4276 (
            .O(N__18854),
            .I(N__18847));
    LocalMux I__4275 (
            .O(N__18847),
            .I(N__18844));
    Odrv4 I__4274 (
            .O(N__18844),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    InMux I__4273 (
            .O(N__18841),
            .I(N__18835));
    InMux I__4272 (
            .O(N__18840),
            .I(N__18835));
    LocalMux I__4271 (
            .O(N__18835),
            .I(N__18832));
    Odrv4 I__4270 (
            .O(N__18832),
            .I(\Lab_UT.dictrl.N_33_0 ));
    InMux I__4269 (
            .O(N__18829),
            .I(N__18826));
    LocalMux I__4268 (
            .O(N__18826),
            .I(N__18823));
    Odrv4 I__4267 (
            .O(N__18823),
            .I(\Lab_UT.dictrl.N_60_0_0 ));
    CascadeMux I__4266 (
            .O(N__18820),
            .I(\Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ));
    InMux I__4265 (
            .O(N__18817),
            .I(N__18805));
    InMux I__4264 (
            .O(N__18816),
            .I(N__18805));
    InMux I__4263 (
            .O(N__18815),
            .I(N__18805));
    InMux I__4262 (
            .O(N__18814),
            .I(N__18805));
    LocalMux I__4261 (
            .O(N__18805),
            .I(\Lab_UT.dictrl.N_26_0 ));
    InMux I__4260 (
            .O(N__18802),
            .I(N__18796));
    InMux I__4259 (
            .O(N__18801),
            .I(N__18796));
    LocalMux I__4258 (
            .O(N__18796),
            .I(N__18793));
    Span4Mux_v I__4257 (
            .O(N__18793),
            .I(N__18790));
    Odrv4 I__4256 (
            .O(N__18790),
            .I(\Lab_UT.dictrl.i8_mux_0 ));
    CascadeMux I__4255 (
            .O(N__18787),
            .I(N__18784));
    InMux I__4254 (
            .O(N__18784),
            .I(N__18781));
    LocalMux I__4253 (
            .O(N__18781),
            .I(\Lab_UT.dictrl.m34_0 ));
    InMux I__4252 (
            .O(N__18778),
            .I(N__18774));
    InMux I__4251 (
            .O(N__18777),
            .I(N__18771));
    LocalMux I__4250 (
            .O(N__18774),
            .I(N__18764));
    LocalMux I__4249 (
            .O(N__18771),
            .I(N__18764));
    CascadeMux I__4248 (
            .O(N__18770),
            .I(N__18761));
    CascadeMux I__4247 (
            .O(N__18769),
            .I(N__18758));
    Span4Mux_h I__4246 (
            .O(N__18764),
            .I(N__18755));
    InMux I__4245 (
            .O(N__18761),
            .I(N__18750));
    InMux I__4244 (
            .O(N__18758),
            .I(N__18750));
    Odrv4 I__4243 (
            .O(N__18755),
            .I(\Lab_UT.dictrl.N_18 ));
    LocalMux I__4242 (
            .O(N__18750),
            .I(\Lab_UT.dictrl.N_18 ));
    CascadeMux I__4241 (
            .O(N__18745),
            .I(N__18742));
    InMux I__4240 (
            .O(N__18742),
            .I(N__18737));
    CascadeMux I__4239 (
            .O(N__18741),
            .I(N__18734));
    CascadeMux I__4238 (
            .O(N__18740),
            .I(N__18730));
    LocalMux I__4237 (
            .O(N__18737),
            .I(N__18727));
    InMux I__4236 (
            .O(N__18734),
            .I(N__18723));
    InMux I__4235 (
            .O(N__18733),
            .I(N__18718));
    InMux I__4234 (
            .O(N__18730),
            .I(N__18718));
    Span4Mux_h I__4233 (
            .O(N__18727),
            .I(N__18715));
    InMux I__4232 (
            .O(N__18726),
            .I(N__18712));
    LocalMux I__4231 (
            .O(N__18723),
            .I(N__18709));
    LocalMux I__4230 (
            .O(N__18718),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    Odrv4 I__4229 (
            .O(N__18715),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    LocalMux I__4228 (
            .O(N__18712),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    Odrv12 I__4227 (
            .O(N__18709),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    CascadeMux I__4226 (
            .O(N__18700),
            .I(N__18696));
    InMux I__4225 (
            .O(N__18699),
            .I(N__18690));
    InMux I__4224 (
            .O(N__18696),
            .I(N__18690));
    InMux I__4223 (
            .O(N__18695),
            .I(N__18687));
    LocalMux I__4222 (
            .O(N__18690),
            .I(N__18684));
    LocalMux I__4221 (
            .O(N__18687),
            .I(N__18681));
    Span4Mux_h I__4220 (
            .O(N__18684),
            .I(N__18678));
    Span4Mux_h I__4219 (
            .O(N__18681),
            .I(N__18675));
    Odrv4 I__4218 (
            .O(N__18678),
            .I(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ));
    Odrv4 I__4217 (
            .O(N__18675),
            .I(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ));
    InMux I__4216 (
            .O(N__18670),
            .I(N__18667));
    LocalMux I__4215 (
            .O(N__18667),
            .I(\Lab_UT.dictrl.g0_1_mb_rn_0 ));
    CascadeMux I__4214 (
            .O(N__18664),
            .I(\Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ));
    InMux I__4213 (
            .O(N__18661),
            .I(N__18658));
    LocalMux I__4212 (
            .O(N__18658),
            .I(N__18654));
    InMux I__4211 (
            .O(N__18657),
            .I(N__18651));
    Span4Mux_h I__4210 (
            .O(N__18654),
            .I(N__18648));
    LocalMux I__4209 (
            .O(N__18651),
            .I(N__18645));
    Span4Mux_v I__4208 (
            .O(N__18648),
            .I(N__18642));
    Span4Mux_h I__4207 (
            .O(N__18645),
            .I(N__18639));
    Odrv4 I__4206 (
            .O(N__18642),
            .I(\Lab_UT.dictrl.N_57_1 ));
    Odrv4 I__4205 (
            .O(N__18639),
            .I(\Lab_UT.dictrl.N_57_1 ));
    CascadeMux I__4204 (
            .O(N__18634),
            .I(N__18631));
    InMux I__4203 (
            .O(N__18631),
            .I(N__18627));
    CascadeMux I__4202 (
            .O(N__18630),
            .I(N__18624));
    LocalMux I__4201 (
            .O(N__18627),
            .I(N__18621));
    InMux I__4200 (
            .O(N__18624),
            .I(N__18618));
    Span4Mux_s3_v I__4199 (
            .O(N__18621),
            .I(N__18615));
    LocalMux I__4198 (
            .O(N__18618),
            .I(N__18612));
    Span4Mux_v I__4197 (
            .O(N__18615),
            .I(N__18607));
    Span4Mux_s3_h I__4196 (
            .O(N__18612),
            .I(N__18607));
    Span4Mux_h I__4195 (
            .O(N__18607),
            .I(N__18604));
    Odrv4 I__4194 (
            .O(N__18604),
            .I(\Lab_UT.dictrl.N_55_1 ));
    CascadeMux I__4193 (
            .O(N__18601),
            .I(N__18598));
    InMux I__4192 (
            .O(N__18598),
            .I(N__18594));
    CascadeMux I__4191 (
            .O(N__18597),
            .I(N__18590));
    LocalMux I__4190 (
            .O(N__18594),
            .I(N__18587));
    InMux I__4189 (
            .O(N__18593),
            .I(N__18582));
    InMux I__4188 (
            .O(N__18590),
            .I(N__18582));
    Span4Mux_v I__4187 (
            .O(N__18587),
            .I(N__18579));
    LocalMux I__4186 (
            .O(N__18582),
            .I(N__18576));
    Span4Mux_v I__4185 (
            .O(N__18579),
            .I(N__18573));
    Span4Mux_v I__4184 (
            .O(N__18576),
            .I(N__18570));
    Odrv4 I__4183 (
            .O(N__18573),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    Odrv4 I__4182 (
            .O(N__18570),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    CascadeMux I__4181 (
            .O(N__18565),
            .I(\Lab_UT.dictrl.next_state_1_2_cascade_ ));
    InMux I__4180 (
            .O(N__18562),
            .I(N__18552));
    InMux I__4179 (
            .O(N__18561),
            .I(N__18552));
    InMux I__4178 (
            .O(N__18560),
            .I(N__18552));
    CascadeMux I__4177 (
            .O(N__18559),
            .I(N__18549));
    LocalMux I__4176 (
            .O(N__18552),
            .I(N__18546));
    InMux I__4175 (
            .O(N__18549),
            .I(N__18543));
    Odrv4 I__4174 (
            .O(N__18546),
            .I(\Lab_UT.dictrl.state_i_4_2 ));
    LocalMux I__4173 (
            .O(N__18543),
            .I(\Lab_UT.dictrl.state_i_4_2 ));
    CEMux I__4172 (
            .O(N__18538),
            .I(N__18534));
    CEMux I__4171 (
            .O(N__18537),
            .I(N__18531));
    LocalMux I__4170 (
            .O(N__18534),
            .I(N__18527));
    LocalMux I__4169 (
            .O(N__18531),
            .I(N__18523));
    CEMux I__4168 (
            .O(N__18530),
            .I(N__18520));
    Span4Mux_h I__4167 (
            .O(N__18527),
            .I(N__18517));
    CEMux I__4166 (
            .O(N__18526),
            .I(N__18514));
    Span4Mux_s3_h I__4165 (
            .O(N__18523),
            .I(N__18509));
    LocalMux I__4164 (
            .O(N__18520),
            .I(N__18509));
    Sp12to4 I__4163 (
            .O(N__18517),
            .I(N__18506));
    LocalMux I__4162 (
            .O(N__18514),
            .I(N__18501));
    Span4Mux_h I__4161 (
            .O(N__18509),
            .I(N__18501));
    Odrv12 I__4160 (
            .O(N__18506),
            .I(\Lab_UT.bu_rx_data_rdy_0 ));
    Odrv4 I__4159 (
            .O(N__18501),
            .I(\Lab_UT.bu_rx_data_rdy_0 ));
    InMux I__4158 (
            .O(N__18496),
            .I(N__18490));
    InMux I__4157 (
            .O(N__18495),
            .I(N__18490));
    LocalMux I__4156 (
            .O(N__18490),
            .I(\Lab_UT.dictrl.g0_1_mb_sn ));
    InMux I__4155 (
            .O(N__18487),
            .I(N__18483));
    InMux I__4154 (
            .O(N__18486),
            .I(N__18479));
    LocalMux I__4153 (
            .O(N__18483),
            .I(N__18476));
    InMux I__4152 (
            .O(N__18482),
            .I(N__18473));
    LocalMux I__4151 (
            .O(N__18479),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    Odrv4 I__4150 (
            .O(N__18476),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    LocalMux I__4149 (
            .O(N__18473),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    CascadeMux I__4148 (
            .O(N__18466),
            .I(\Lab_UT.dictrl.un15_loadalarm_0_cascade_ ));
    InMux I__4147 (
            .O(N__18463),
            .I(N__18460));
    LocalMux I__4146 (
            .O(N__18460),
            .I(\Lab_UT.dictrl.loadalarm_0_0 ));
    InMux I__4145 (
            .O(N__18457),
            .I(N__18452));
    CascadeMux I__4144 (
            .O(N__18456),
            .I(N__18449));
    CascadeMux I__4143 (
            .O(N__18455),
            .I(N__18444));
    LocalMux I__4142 (
            .O(N__18452),
            .I(N__18441));
    InMux I__4141 (
            .O(N__18449),
            .I(N__18438));
    CascadeMux I__4140 (
            .O(N__18448),
            .I(N__18435));
    InMux I__4139 (
            .O(N__18447),
            .I(N__18429));
    InMux I__4138 (
            .O(N__18444),
            .I(N__18423));
    Span4Mux_v I__4137 (
            .O(N__18441),
            .I(N__18418));
    LocalMux I__4136 (
            .O(N__18438),
            .I(N__18418));
    InMux I__4135 (
            .O(N__18435),
            .I(N__18412));
    InMux I__4134 (
            .O(N__18434),
            .I(N__18405));
    InMux I__4133 (
            .O(N__18433),
            .I(N__18405));
    InMux I__4132 (
            .O(N__18432),
            .I(N__18405));
    LocalMux I__4131 (
            .O(N__18429),
            .I(N__18402));
    InMux I__4130 (
            .O(N__18428),
            .I(N__18395));
    InMux I__4129 (
            .O(N__18427),
            .I(N__18395));
    InMux I__4128 (
            .O(N__18426),
            .I(N__18395));
    LocalMux I__4127 (
            .O(N__18423),
            .I(N__18390));
    Span4Mux_h I__4126 (
            .O(N__18418),
            .I(N__18390));
    InMux I__4125 (
            .O(N__18417),
            .I(N__18383));
    InMux I__4124 (
            .O(N__18416),
            .I(N__18383));
    InMux I__4123 (
            .O(N__18415),
            .I(N__18383));
    LocalMux I__4122 (
            .O(N__18412),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4121 (
            .O(N__18405),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__4120 (
            .O(N__18402),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4119 (
            .O(N__18395),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__4118 (
            .O(N__18390),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4117 (
            .O(N__18383),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    InMux I__4116 (
            .O(N__18370),
            .I(N__18365));
    InMux I__4115 (
            .O(N__18369),
            .I(N__18351));
    InMux I__4114 (
            .O(N__18368),
            .I(N__18351));
    LocalMux I__4113 (
            .O(N__18365),
            .I(N__18346));
    InMux I__4112 (
            .O(N__18364),
            .I(N__18341));
    InMux I__4111 (
            .O(N__18363),
            .I(N__18341));
    InMux I__4110 (
            .O(N__18362),
            .I(N__18332));
    InMux I__4109 (
            .O(N__18361),
            .I(N__18332));
    InMux I__4108 (
            .O(N__18360),
            .I(N__18332));
    InMux I__4107 (
            .O(N__18359),
            .I(N__18332));
    InMux I__4106 (
            .O(N__18358),
            .I(N__18327));
    InMux I__4105 (
            .O(N__18357),
            .I(N__18327));
    InMux I__4104 (
            .O(N__18356),
            .I(N__18321));
    LocalMux I__4103 (
            .O(N__18351),
            .I(N__18316));
    InMux I__4102 (
            .O(N__18350),
            .I(N__18311));
    InMux I__4101 (
            .O(N__18349),
            .I(N__18311));
    Span4Mux_v I__4100 (
            .O(N__18346),
            .I(N__18308));
    LocalMux I__4099 (
            .O(N__18341),
            .I(N__18301));
    LocalMux I__4098 (
            .O(N__18332),
            .I(N__18301));
    LocalMux I__4097 (
            .O(N__18327),
            .I(N__18301));
    InMux I__4096 (
            .O(N__18326),
            .I(N__18294));
    InMux I__4095 (
            .O(N__18325),
            .I(N__18294));
    InMux I__4094 (
            .O(N__18324),
            .I(N__18294));
    LocalMux I__4093 (
            .O(N__18321),
            .I(N__18291));
    InMux I__4092 (
            .O(N__18320),
            .I(N__18286));
    InMux I__4091 (
            .O(N__18319),
            .I(N__18286));
    Span4Mux_v I__4090 (
            .O(N__18316),
            .I(N__18283));
    LocalMux I__4089 (
            .O(N__18311),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__4088 (
            .O(N__18308),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__4087 (
            .O(N__18301),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__4086 (
            .O(N__18294),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__4085 (
            .O(N__18291),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__4084 (
            .O(N__18286),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__4083 (
            .O(N__18283),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    CascadeMux I__4082 (
            .O(N__18268),
            .I(N__18262));
    InMux I__4081 (
            .O(N__18267),
            .I(N__18253));
    InMux I__4080 (
            .O(N__18266),
            .I(N__18253));
    InMux I__4079 (
            .O(N__18265),
            .I(N__18253));
    InMux I__4078 (
            .O(N__18262),
            .I(N__18249));
    CascadeMux I__4077 (
            .O(N__18261),
            .I(N__18245));
    InMux I__4076 (
            .O(N__18260),
            .I(N__18239));
    LocalMux I__4075 (
            .O(N__18253),
            .I(N__18236));
    InMux I__4074 (
            .O(N__18252),
            .I(N__18233));
    LocalMux I__4073 (
            .O(N__18249),
            .I(N__18230));
    InMux I__4072 (
            .O(N__18248),
            .I(N__18227));
    InMux I__4071 (
            .O(N__18245),
            .I(N__18222));
    InMux I__4070 (
            .O(N__18244),
            .I(N__18222));
    InMux I__4069 (
            .O(N__18243),
            .I(N__18217));
    InMux I__4068 (
            .O(N__18242),
            .I(N__18217));
    LocalMux I__4067 (
            .O(N__18239),
            .I(N__18213));
    Span4Mux_h I__4066 (
            .O(N__18236),
            .I(N__18208));
    LocalMux I__4065 (
            .O(N__18233),
            .I(N__18208));
    Span4Mux_v I__4064 (
            .O(N__18230),
            .I(N__18203));
    LocalMux I__4063 (
            .O(N__18227),
            .I(N__18203));
    LocalMux I__4062 (
            .O(N__18222),
            .I(N__18198));
    LocalMux I__4061 (
            .O(N__18217),
            .I(N__18198));
    InMux I__4060 (
            .O(N__18216),
            .I(N__18195));
    Span4Mux_h I__4059 (
            .O(N__18213),
            .I(N__18192));
    Span4Mux_h I__4058 (
            .O(N__18208),
            .I(N__18189));
    Span4Mux_h I__4057 (
            .O(N__18203),
            .I(N__18186));
    Span12Mux_s8_h I__4056 (
            .O(N__18198),
            .I(N__18183));
    LocalMux I__4055 (
            .O(N__18195),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__4054 (
            .O(N__18192),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__4053 (
            .O(N__18189),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__4052 (
            .O(N__18186),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv12 I__4051 (
            .O(N__18183),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    InMux I__4050 (
            .O(N__18172),
            .I(N__18160));
    InMux I__4049 (
            .O(N__18171),
            .I(N__18160));
    InMux I__4048 (
            .O(N__18170),
            .I(N__18160));
    InMux I__4047 (
            .O(N__18169),
            .I(N__18160));
    LocalMux I__4046 (
            .O(N__18160),
            .I(N__18154));
    InMux I__4045 (
            .O(N__18159),
            .I(N__18150));
    InMux I__4044 (
            .O(N__18158),
            .I(N__18147));
    InMux I__4043 (
            .O(N__18157),
            .I(N__18144));
    Span4Mux_s3_h I__4042 (
            .O(N__18154),
            .I(N__18141));
    InMux I__4041 (
            .O(N__18153),
            .I(N__18138));
    LocalMux I__4040 (
            .O(N__18150),
            .I(N__18133));
    LocalMux I__4039 (
            .O(N__18147),
            .I(N__18133));
    LocalMux I__4038 (
            .O(N__18144),
            .I(\Lab_UT.next_state_1 ));
    Odrv4 I__4037 (
            .O(N__18141),
            .I(\Lab_UT.next_state_1 ));
    LocalMux I__4036 (
            .O(N__18138),
            .I(\Lab_UT.next_state_1 ));
    Odrv12 I__4035 (
            .O(N__18133),
            .I(\Lab_UT.next_state_1 ));
    InMux I__4034 (
            .O(N__18124),
            .I(N__18115));
    InMux I__4033 (
            .O(N__18123),
            .I(N__18106));
    InMux I__4032 (
            .O(N__18122),
            .I(N__18106));
    InMux I__4031 (
            .O(N__18121),
            .I(N__18106));
    InMux I__4030 (
            .O(N__18120),
            .I(N__18106));
    InMux I__4029 (
            .O(N__18119),
            .I(N__18103));
    InMux I__4028 (
            .O(N__18118),
            .I(N__18100));
    LocalMux I__4027 (
            .O(N__18115),
            .I(N__18097));
    LocalMux I__4026 (
            .O(N__18106),
            .I(\Lab_UT.next_state_2 ));
    LocalMux I__4025 (
            .O(N__18103),
            .I(\Lab_UT.next_state_2 ));
    LocalMux I__4024 (
            .O(N__18100),
            .I(\Lab_UT.next_state_2 ));
    Odrv4 I__4023 (
            .O(N__18097),
            .I(\Lab_UT.next_state_2 ));
    CascadeMux I__4022 (
            .O(N__18088),
            .I(N__18084));
    CascadeMux I__4021 (
            .O(N__18087),
            .I(N__18080));
    InMux I__4020 (
            .O(N__18084),
            .I(N__18075));
    InMux I__4019 (
            .O(N__18083),
            .I(N__18068));
    InMux I__4018 (
            .O(N__18080),
            .I(N__18068));
    InMux I__4017 (
            .O(N__18079),
            .I(N__18068));
    InMux I__4016 (
            .O(N__18078),
            .I(N__18062));
    LocalMux I__4015 (
            .O(N__18075),
            .I(N__18057));
    LocalMux I__4014 (
            .O(N__18068),
            .I(N__18057));
    InMux I__4013 (
            .O(N__18067),
            .I(N__18050));
    InMux I__4012 (
            .O(N__18066),
            .I(N__18050));
    InMux I__4011 (
            .O(N__18065),
            .I(N__18050));
    LocalMux I__4010 (
            .O(N__18062),
            .I(N__18047));
    Span4Mux_v I__4009 (
            .O(N__18057),
            .I(N__18041));
    LocalMux I__4008 (
            .O(N__18050),
            .I(N__18041));
    Span4Mux_v I__4007 (
            .O(N__18047),
            .I(N__18037));
    InMux I__4006 (
            .O(N__18046),
            .I(N__18034));
    Span4Mux_h I__4005 (
            .O(N__18041),
            .I(N__18031));
    InMux I__4004 (
            .O(N__18040),
            .I(N__18028));
    Sp12to4 I__4003 (
            .O(N__18037),
            .I(N__18023));
    LocalMux I__4002 (
            .O(N__18034),
            .I(N__18023));
    Span4Mux_h I__4001 (
            .O(N__18031),
            .I(N__18020));
    LocalMux I__4000 (
            .O(N__18028),
            .I(bu_rx_data_rdy));
    Odrv12 I__3999 (
            .O(N__18023),
            .I(bu_rx_data_rdy));
    Odrv4 I__3998 (
            .O(N__18020),
            .I(bu_rx_data_rdy));
    CascadeMux I__3997 (
            .O(N__18013),
            .I(N__18008));
    InMux I__3996 (
            .O(N__18012),
            .I(N__18005));
    CascadeMux I__3995 (
            .O(N__18011),
            .I(N__18002));
    InMux I__3994 (
            .O(N__18008),
            .I(N__17999));
    LocalMux I__3993 (
            .O(N__18005),
            .I(N__17996));
    InMux I__3992 (
            .O(N__18002),
            .I(N__17993));
    LocalMux I__3991 (
            .O(N__17999),
            .I(N__17989));
    Span4Mux_v I__3990 (
            .O(N__17996),
            .I(N__17984));
    LocalMux I__3989 (
            .O(N__17993),
            .I(N__17984));
    InMux I__3988 (
            .O(N__17992),
            .I(N__17981));
    Span4Mux_v I__3987 (
            .O(N__17989),
            .I(N__17978));
    Odrv4 I__3986 (
            .O(N__17984),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    LocalMux I__3985 (
            .O(N__17981),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    Odrv4 I__3984 (
            .O(N__17978),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    CascadeMux I__3983 (
            .O(N__17971),
            .I(\Lab_UT.didp.countrce3.q_5_1_cascade_ ));
    InMux I__3982 (
            .O(N__17968),
            .I(N__17965));
    LocalMux I__3981 (
            .O(N__17965),
            .I(N__17961));
    InMux I__3980 (
            .O(N__17964),
            .I(N__17958));
    Span4Mux_v I__3979 (
            .O(N__17961),
            .I(N__17953));
    LocalMux I__3978 (
            .O(N__17958),
            .I(N__17953));
    Span4Mux_h I__3977 (
            .O(N__17953),
            .I(N__17949));
    InMux I__3976 (
            .O(N__17952),
            .I(N__17946));
    Odrv4 I__3975 (
            .O(N__17949),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    LocalMux I__3974 (
            .O(N__17946),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    InMux I__3973 (
            .O(N__17941),
            .I(N__17937));
    CascadeMux I__3972 (
            .O(N__17940),
            .I(N__17934));
    LocalMux I__3971 (
            .O(N__17937),
            .I(N__17926));
    InMux I__3970 (
            .O(N__17934),
            .I(N__17923));
    InMux I__3969 (
            .O(N__17933),
            .I(N__17920));
    InMux I__3968 (
            .O(N__17932),
            .I(N__17913));
    InMux I__3967 (
            .O(N__17931),
            .I(N__17913));
    InMux I__3966 (
            .O(N__17930),
            .I(N__17913));
    InMux I__3965 (
            .O(N__17929),
            .I(N__17910));
    Span4Mux_v I__3964 (
            .O(N__17926),
            .I(N__17905));
    LocalMux I__3963 (
            .O(N__17923),
            .I(N__17905));
    LocalMux I__3962 (
            .O(N__17920),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3961 (
            .O(N__17913),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3960 (
            .O(N__17910),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv4 I__3959 (
            .O(N__17905),
            .I(\Lab_UT.di_Mones_1 ));
    CascadeMux I__3958 (
            .O(N__17896),
            .I(N__17891));
    CascadeMux I__3957 (
            .O(N__17895),
            .I(N__17886));
    InMux I__3956 (
            .O(N__17894),
            .I(N__17881));
    InMux I__3955 (
            .O(N__17891),
            .I(N__17881));
    InMux I__3954 (
            .O(N__17890),
            .I(N__17878));
    InMux I__3953 (
            .O(N__17889),
            .I(N__17873));
    InMux I__3952 (
            .O(N__17886),
            .I(N__17873));
    LocalMux I__3951 (
            .O(N__17881),
            .I(N__17870));
    LocalMux I__3950 (
            .O(N__17878),
            .I(N__17866));
    LocalMux I__3949 (
            .O(N__17873),
            .I(N__17863));
    Span4Mux_v I__3948 (
            .O(N__17870),
            .I(N__17860));
    InMux I__3947 (
            .O(N__17869),
            .I(N__17857));
    Span4Mux_v I__3946 (
            .O(N__17866),
            .I(N__17854));
    Span12Mux_s8_h I__3945 (
            .O(N__17863),
            .I(N__17851));
    Span4Mux_h I__3944 (
            .O(N__17860),
            .I(N__17848));
    LocalMux I__3943 (
            .O(N__17857),
            .I(N__17843));
    Span4Mux_s2_v I__3942 (
            .O(N__17854),
            .I(N__17843));
    Odrv12 I__3941 (
            .O(N__17851),
            .I(\Lab_UT.state_ret_8_ess ));
    Odrv4 I__3940 (
            .O(N__17848),
            .I(\Lab_UT.state_ret_8_ess ));
    Odrv4 I__3939 (
            .O(N__17843),
            .I(\Lab_UT.state_ret_8_ess ));
    CascadeMux I__3938 (
            .O(N__17836),
            .I(N__17832));
    CascadeMux I__3937 (
            .O(N__17835),
            .I(N__17828));
    InMux I__3936 (
            .O(N__17832),
            .I(N__17815));
    InMux I__3935 (
            .O(N__17831),
            .I(N__17815));
    InMux I__3934 (
            .O(N__17828),
            .I(N__17815));
    InMux I__3933 (
            .O(N__17827),
            .I(N__17815));
    InMux I__3932 (
            .O(N__17826),
            .I(N__17810));
    InMux I__3931 (
            .O(N__17825),
            .I(N__17810));
    InMux I__3930 (
            .O(N__17824),
            .I(N__17806));
    LocalMux I__3929 (
            .O(N__17815),
            .I(N__17803));
    LocalMux I__3928 (
            .O(N__17810),
            .I(N__17800));
    InMux I__3927 (
            .O(N__17809),
            .I(N__17797));
    LocalMux I__3926 (
            .O(N__17806),
            .I(\Lab_UT.next_state_0 ));
    Odrv4 I__3925 (
            .O(N__17803),
            .I(\Lab_UT.next_state_0 ));
    Odrv12 I__3924 (
            .O(N__17800),
            .I(\Lab_UT.next_state_0 ));
    LocalMux I__3923 (
            .O(N__17797),
            .I(\Lab_UT.next_state_0 ));
    InMux I__3922 (
            .O(N__17788),
            .I(N__17785));
    LocalMux I__3921 (
            .O(N__17785),
            .I(N__17782));
    Odrv12 I__3920 (
            .O(N__17782),
            .I(\Lab_UT.didp.N_90 ));
    InMux I__3919 (
            .O(N__17779),
            .I(N__17776));
    LocalMux I__3918 (
            .O(N__17776),
            .I(N__17773));
    Odrv12 I__3917 (
            .O(N__17773),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__3916 (
            .O(N__17770),
            .I(N__17767));
    LocalMux I__3915 (
            .O(N__17767),
            .I(\Lab_UT.LdSones_i_4 ));
    CascadeMux I__3914 (
            .O(N__17764),
            .I(N__17759));
    InMux I__3913 (
            .O(N__17763),
            .I(N__17756));
    InMux I__3912 (
            .O(N__17762),
            .I(N__17753));
    InMux I__3911 (
            .O(N__17759),
            .I(N__17750));
    LocalMux I__3910 (
            .O(N__17756),
            .I(N__17747));
    LocalMux I__3909 (
            .O(N__17753),
            .I(N__17739));
    LocalMux I__3908 (
            .O(N__17750),
            .I(N__17739));
    Span4Mux_h I__3907 (
            .O(N__17747),
            .I(N__17739));
    InMux I__3906 (
            .O(N__17746),
            .I(N__17736));
    Span4Mux_h I__3905 (
            .O(N__17739),
            .I(N__17733));
    LocalMux I__3904 (
            .O(N__17736),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    Odrv4 I__3903 (
            .O(N__17733),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    InMux I__3902 (
            .O(N__17728),
            .I(N__17722));
    InMux I__3901 (
            .O(N__17727),
            .I(N__17718));
    InMux I__3900 (
            .O(N__17726),
            .I(N__17714));
    InMux I__3899 (
            .O(N__17725),
            .I(N__17711));
    LocalMux I__3898 (
            .O(N__17722),
            .I(N__17708));
    InMux I__3897 (
            .O(N__17721),
            .I(N__17705));
    LocalMux I__3896 (
            .O(N__17718),
            .I(N__17702));
    InMux I__3895 (
            .O(N__17717),
            .I(N__17699));
    LocalMux I__3894 (
            .O(N__17714),
            .I(N__17696));
    LocalMux I__3893 (
            .O(N__17711),
            .I(N__17693));
    Span4Mux_h I__3892 (
            .O(N__17708),
            .I(N__17690));
    LocalMux I__3891 (
            .O(N__17705),
            .I(N__17681));
    Span4Mux_h I__3890 (
            .O(N__17702),
            .I(N__17681));
    LocalMux I__3889 (
            .O(N__17699),
            .I(N__17681));
    Span4Mux_h I__3888 (
            .O(N__17696),
            .I(N__17678));
    Span4Mux_s2_v I__3887 (
            .O(N__17693),
            .I(N__17675));
    Span4Mux_v I__3886 (
            .O(N__17690),
            .I(N__17672));
    InMux I__3885 (
            .O(N__17689),
            .I(N__17667));
    InMux I__3884 (
            .O(N__17688),
            .I(N__17667));
    Span4Mux_h I__3883 (
            .O(N__17681),
            .I(N__17664));
    Span4Mux_h I__3882 (
            .O(N__17678),
            .I(N__17659));
    Span4Mux_h I__3881 (
            .O(N__17675),
            .I(N__17659));
    Odrv4 I__3880 (
            .O(N__17672),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3879 (
            .O(N__17667),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__3878 (
            .O(N__17664),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__3877 (
            .O(N__17659),
            .I(\Lab_UT.di_Sones_0 ));
    InMux I__3876 (
            .O(N__17650),
            .I(N__17647));
    LocalMux I__3875 (
            .O(N__17647),
            .I(N__17643));
    InMux I__3874 (
            .O(N__17646),
            .I(N__17640));
    Span4Mux_v I__3873 (
            .O(N__17643),
            .I(N__17635));
    LocalMux I__3872 (
            .O(N__17640),
            .I(N__17632));
    InMux I__3871 (
            .O(N__17639),
            .I(N__17629));
    CascadeMux I__3870 (
            .O(N__17638),
            .I(N__17626));
    Span4Mux_h I__3869 (
            .O(N__17635),
            .I(N__17623));
    Span4Mux_v I__3868 (
            .O(N__17632),
            .I(N__17620));
    LocalMux I__3867 (
            .O(N__17629),
            .I(N__17617));
    InMux I__3866 (
            .O(N__17626),
            .I(N__17614));
    Odrv4 I__3865 (
            .O(N__17623),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__3864 (
            .O(N__17620),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__3863 (
            .O(N__17617),
            .I(\Lab_UT.LdSones ));
    LocalMux I__3862 (
            .O(N__17614),
            .I(\Lab_UT.LdSones ));
    InMux I__3861 (
            .O(N__17605),
            .I(N__17595));
    InMux I__3860 (
            .O(N__17604),
            .I(N__17595));
    InMux I__3859 (
            .O(N__17603),
            .I(N__17595));
    InMux I__3858 (
            .O(N__17602),
            .I(N__17592));
    LocalMux I__3857 (
            .O(N__17595),
            .I(N__17586));
    LocalMux I__3856 (
            .O(N__17592),
            .I(N__17583));
    InMux I__3855 (
            .O(N__17591),
            .I(N__17579));
    InMux I__3854 (
            .O(N__17590),
            .I(N__17575));
    InMux I__3853 (
            .O(N__17589),
            .I(N__17572));
    Span4Mux_h I__3852 (
            .O(N__17586),
            .I(N__17569));
    Span4Mux_h I__3851 (
            .O(N__17583),
            .I(N__17566));
    InMux I__3850 (
            .O(N__17582),
            .I(N__17563));
    LocalMux I__3849 (
            .O(N__17579),
            .I(N__17560));
    InMux I__3848 (
            .O(N__17578),
            .I(N__17557));
    LocalMux I__3847 (
            .O(N__17575),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3846 (
            .O(N__17572),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3845 (
            .O(N__17569),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3844 (
            .O(N__17566),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3843 (
            .O(N__17563),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3842 (
            .O(N__17560),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3841 (
            .O(N__17557),
            .I(\Lab_UT.di_Sones_1 ));
    InMux I__3840 (
            .O(N__17542),
            .I(N__17539));
    LocalMux I__3839 (
            .O(N__17539),
            .I(N__17536));
    Odrv4 I__3838 (
            .O(N__17536),
            .I(\Lab_UT.didp.countrce1.q_5_1 ));
    CascadeMux I__3837 (
            .O(N__17533),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    InMux I__3836 (
            .O(N__17530),
            .I(N__17527));
    LocalMux I__3835 (
            .O(N__17527),
            .I(\Lab_UT.didp.countrce3.q_5_3 ));
    CascadeMux I__3834 (
            .O(N__17524),
            .I(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ));
    InMux I__3833 (
            .O(N__17521),
            .I(N__17511));
    InMux I__3832 (
            .O(N__17520),
            .I(N__17511));
    InMux I__3831 (
            .O(N__17519),
            .I(N__17511));
    InMux I__3830 (
            .O(N__17518),
            .I(N__17496));
    LocalMux I__3829 (
            .O(N__17511),
            .I(N__17493));
    InMux I__3828 (
            .O(N__17510),
            .I(N__17490));
    InMux I__3827 (
            .O(N__17509),
            .I(N__17479));
    InMux I__3826 (
            .O(N__17508),
            .I(N__17479));
    InMux I__3825 (
            .O(N__17507),
            .I(N__17479));
    InMux I__3824 (
            .O(N__17506),
            .I(N__17479));
    InMux I__3823 (
            .O(N__17505),
            .I(N__17479));
    InMux I__3822 (
            .O(N__17504),
            .I(N__17470));
    InMux I__3821 (
            .O(N__17503),
            .I(N__17470));
    InMux I__3820 (
            .O(N__17502),
            .I(N__17470));
    InMux I__3819 (
            .O(N__17501),
            .I(N__17470));
    InMux I__3818 (
            .O(N__17500),
            .I(N__17467));
    InMux I__3817 (
            .O(N__17499),
            .I(N__17464));
    LocalMux I__3816 (
            .O(N__17496),
            .I(N__17461));
    Span4Mux_h I__3815 (
            .O(N__17493),
            .I(N__17456));
    LocalMux I__3814 (
            .O(N__17490),
            .I(N__17456));
    LocalMux I__3813 (
            .O(N__17479),
            .I(N__17451));
    LocalMux I__3812 (
            .O(N__17470),
            .I(N__17451));
    LocalMux I__3811 (
            .O(N__17467),
            .I(\Lab_UT.loadalarm_0 ));
    LocalMux I__3810 (
            .O(N__17464),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv4 I__3809 (
            .O(N__17461),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv4 I__3808 (
            .O(N__17456),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv12 I__3807 (
            .O(N__17451),
            .I(\Lab_UT.loadalarm_0 ));
    InMux I__3806 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__3805 (
            .O(N__17437),
            .I(N__17434));
    Span4Mux_h I__3804 (
            .O(N__17434),
            .I(N__17426));
    InMux I__3803 (
            .O(N__17433),
            .I(N__17423));
    InMux I__3802 (
            .O(N__17432),
            .I(N__17418));
    InMux I__3801 (
            .O(N__17431),
            .I(N__17418));
    InMux I__3800 (
            .O(N__17430),
            .I(N__17415));
    InMux I__3799 (
            .O(N__17429),
            .I(N__17412));
    Odrv4 I__3798 (
            .O(N__17426),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3797 (
            .O(N__17423),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3796 (
            .O(N__17418),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3795 (
            .O(N__17415),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3794 (
            .O(N__17412),
            .I(\Lab_UT.di_Mtens_2 ));
    InMux I__3793 (
            .O(N__17401),
            .I(N__17398));
    LocalMux I__3792 (
            .O(N__17398),
            .I(N__17393));
    InMux I__3791 (
            .O(N__17397),
            .I(N__17390));
    InMux I__3790 (
            .O(N__17396),
            .I(N__17387));
    Span4Mux_h I__3789 (
            .O(N__17393),
            .I(N__17384));
    LocalMux I__3788 (
            .O(N__17390),
            .I(N__17381));
    LocalMux I__3787 (
            .O(N__17387),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__3786 (
            .O(N__17384),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv12 I__3785 (
            .O(N__17381),
            .I(\Lab_UT.di_AMtens_2 ));
    InMux I__3784 (
            .O(N__17374),
            .I(N__17368));
    CascadeMux I__3783 (
            .O(N__17373),
            .I(N__17364));
    CascadeMux I__3782 (
            .O(N__17372),
            .I(N__17360));
    CascadeMux I__3781 (
            .O(N__17371),
            .I(N__17356));
    LocalMux I__3780 (
            .O(N__17368),
            .I(N__17353));
    InMux I__3779 (
            .O(N__17367),
            .I(N__17340));
    InMux I__3778 (
            .O(N__17364),
            .I(N__17340));
    InMux I__3777 (
            .O(N__17363),
            .I(N__17340));
    InMux I__3776 (
            .O(N__17360),
            .I(N__17340));
    InMux I__3775 (
            .O(N__17359),
            .I(N__17340));
    InMux I__3774 (
            .O(N__17356),
            .I(N__17340));
    Span4Mux_h I__3773 (
            .O(N__17353),
            .I(N__17337));
    LocalMux I__3772 (
            .O(N__17340),
            .I(N__17334));
    Odrv4 I__3771 (
            .O(N__17337),
            .I(\Lab_UT.min1_2 ));
    Odrv12 I__3770 (
            .O(N__17334),
            .I(\Lab_UT.min1_2 ));
    InMux I__3769 (
            .O(N__17329),
            .I(N__17326));
    LocalMux I__3768 (
            .O(N__17326),
            .I(\Lab_UT.didp.countrce1.q_5_2 ));
    CascadeMux I__3767 (
            .O(N__17323),
            .I(N__17320));
    InMux I__3766 (
            .O(N__17320),
            .I(N__17316));
    CascadeMux I__3765 (
            .O(N__17319),
            .I(N__17313));
    LocalMux I__3764 (
            .O(N__17316),
            .I(N__17309));
    InMux I__3763 (
            .O(N__17313),
            .I(N__17306));
    InMux I__3762 (
            .O(N__17312),
            .I(N__17303));
    Sp12to4 I__3761 (
            .O(N__17309),
            .I(N__17297));
    LocalMux I__3760 (
            .O(N__17306),
            .I(N__17297));
    LocalMux I__3759 (
            .O(N__17303),
            .I(N__17294));
    InMux I__3758 (
            .O(N__17302),
            .I(N__17291));
    Span12Mux_s6_h I__3757 (
            .O(N__17297),
            .I(N__17286));
    Span12Mux_s5_h I__3756 (
            .O(N__17294),
            .I(N__17286));
    LocalMux I__3755 (
            .O(N__17291),
            .I(N__17283));
    Odrv12 I__3754 (
            .O(N__17286),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    Odrv4 I__3753 (
            .O(N__17283),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    InMux I__3752 (
            .O(N__17278),
            .I(N__17272));
    InMux I__3751 (
            .O(N__17277),
            .I(N__17272));
    LocalMux I__3750 (
            .O(N__17272),
            .I(N__17266));
    InMux I__3749 (
            .O(N__17271),
            .I(N__17263));
    InMux I__3748 (
            .O(N__17270),
            .I(N__17259));
    InMux I__3747 (
            .O(N__17269),
            .I(N__17256));
    Span4Mux_h I__3746 (
            .O(N__17266),
            .I(N__17253));
    LocalMux I__3745 (
            .O(N__17263),
            .I(N__17250));
    InMux I__3744 (
            .O(N__17262),
            .I(N__17247));
    LocalMux I__3743 (
            .O(N__17259),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3742 (
            .O(N__17256),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__3741 (
            .O(N__17253),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__3740 (
            .O(N__17250),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3739 (
            .O(N__17247),
            .I(\Lab_UT.di_Sones_2 ));
    InMux I__3738 (
            .O(N__17236),
            .I(N__17232));
    InMux I__3737 (
            .O(N__17235),
            .I(N__17228));
    LocalMux I__3736 (
            .O(N__17232),
            .I(N__17222));
    InMux I__3735 (
            .O(N__17231),
            .I(N__17219));
    LocalMux I__3734 (
            .O(N__17228),
            .I(N__17216));
    InMux I__3733 (
            .O(N__17227),
            .I(N__17213));
    InMux I__3732 (
            .O(N__17226),
            .I(N__17208));
    InMux I__3731 (
            .O(N__17225),
            .I(N__17208));
    Span4Mux_h I__3730 (
            .O(N__17222),
            .I(N__17205));
    LocalMux I__3729 (
            .O(N__17219),
            .I(N__17202));
    Span4Mux_h I__3728 (
            .O(N__17216),
            .I(N__17197));
    LocalMux I__3727 (
            .O(N__17213),
            .I(N__17197));
    LocalMux I__3726 (
            .O(N__17208),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3725 (
            .O(N__17205),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv12 I__3724 (
            .O(N__17202),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3723 (
            .O(N__17197),
            .I(\Lab_UT.di_Mones_2 ));
    InMux I__3722 (
            .O(N__17188),
            .I(N__17184));
    CascadeMux I__3721 (
            .O(N__17187),
            .I(N__17181));
    LocalMux I__3720 (
            .O(N__17184),
            .I(N__17177));
    InMux I__3719 (
            .O(N__17181),
            .I(N__17172));
    CascadeMux I__3718 (
            .O(N__17180),
            .I(N__17169));
    Span4Mux_v I__3717 (
            .O(N__17177),
            .I(N__17166));
    InMux I__3716 (
            .O(N__17176),
            .I(N__17163));
    InMux I__3715 (
            .O(N__17175),
            .I(N__17160));
    LocalMux I__3714 (
            .O(N__17172),
            .I(N__17157));
    InMux I__3713 (
            .O(N__17169),
            .I(N__17154));
    Odrv4 I__3712 (
            .O(N__17166),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3711 (
            .O(N__17163),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3710 (
            .O(N__17160),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__3709 (
            .O(N__17157),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3708 (
            .O(N__17154),
            .I(\Lab_UT.di_Mones_3 ));
    InMux I__3707 (
            .O(N__17143),
            .I(N__17134));
    InMux I__3706 (
            .O(N__17142),
            .I(N__17134));
    InMux I__3705 (
            .O(N__17141),
            .I(N__17134));
    LocalMux I__3704 (
            .O(N__17134),
            .I(N__17131));
    Span4Mux_h I__3703 (
            .O(N__17131),
            .I(N__17128));
    Odrv4 I__3702 (
            .O(N__17128),
            .I(\Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ));
    CascadeMux I__3701 (
            .O(N__17125),
            .I(N__17122));
    InMux I__3700 (
            .O(N__17122),
            .I(N__17118));
    InMux I__3699 (
            .O(N__17121),
            .I(N__17114));
    LocalMux I__3698 (
            .O(N__17118),
            .I(N__17111));
    InMux I__3697 (
            .O(N__17117),
            .I(N__17105));
    LocalMux I__3696 (
            .O(N__17114),
            .I(N__17102));
    Span4Mux_v I__3695 (
            .O(N__17111),
            .I(N__17099));
    InMux I__3694 (
            .O(N__17110),
            .I(N__17094));
    InMux I__3693 (
            .O(N__17109),
            .I(N__17094));
    InMux I__3692 (
            .O(N__17108),
            .I(N__17091));
    LocalMux I__3691 (
            .O(N__17105),
            .I(N__17088));
    Sp12to4 I__3690 (
            .O(N__17102),
            .I(N__17081));
    Sp12to4 I__3689 (
            .O(N__17099),
            .I(N__17081));
    LocalMux I__3688 (
            .O(N__17094),
            .I(N__17081));
    LocalMux I__3687 (
            .O(N__17091),
            .I(N__17078));
    Span4Mux_v I__3686 (
            .O(N__17088),
            .I(N__17075));
    Span12Mux_s5_h I__3685 (
            .O(N__17081),
            .I(N__17072));
    Span12Mux_v I__3684 (
            .O(N__17078),
            .I(N__17069));
    Span4Mux_v I__3683 (
            .O(N__17075),
            .I(N__17066));
    Odrv12 I__3682 (
            .O(N__17072),
            .I(\Lab_UT.LdMtens ));
    Odrv12 I__3681 (
            .O(N__17069),
            .I(\Lab_UT.LdMtens ));
    Odrv4 I__3680 (
            .O(N__17066),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__3679 (
            .O(N__17059),
            .I(N__17056));
    InMux I__3678 (
            .O(N__17056),
            .I(N__17053));
    LocalMux I__3677 (
            .O(N__17053),
            .I(\Lab_UT.didp.countrce4.un20_qPone ));
    InMux I__3676 (
            .O(N__17050),
            .I(N__17047));
    LocalMux I__3675 (
            .O(N__17047),
            .I(N__17041));
    InMux I__3674 (
            .O(N__17046),
            .I(N__17037));
    InMux I__3673 (
            .O(N__17045),
            .I(N__17034));
    InMux I__3672 (
            .O(N__17044),
            .I(N__17031));
    Span4Mux_h I__3671 (
            .O(N__17041),
            .I(N__17028));
    InMux I__3670 (
            .O(N__17040),
            .I(N__17025));
    LocalMux I__3669 (
            .O(N__17037),
            .I(N__17022));
    LocalMux I__3668 (
            .O(N__17034),
            .I(N__17019));
    LocalMux I__3667 (
            .O(N__17031),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__3666 (
            .O(N__17028),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__3665 (
            .O(N__17025),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__3664 (
            .O(N__17022),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__3663 (
            .O(N__17019),
            .I(\Lab_UT.di_Mtens_3 ));
    InMux I__3662 (
            .O(N__17008),
            .I(N__17005));
    LocalMux I__3661 (
            .O(N__17005),
            .I(\Lab_UT.didp.countrce4.q_5_3 ));
    InMux I__3660 (
            .O(N__17002),
            .I(N__16997));
    InMux I__3659 (
            .O(N__17001),
            .I(N__16989));
    InMux I__3658 (
            .O(N__17000),
            .I(N__16989));
    LocalMux I__3657 (
            .O(N__16997),
            .I(N__16986));
    InMux I__3656 (
            .O(N__16996),
            .I(N__16982));
    InMux I__3655 (
            .O(N__16995),
            .I(N__16977));
    InMux I__3654 (
            .O(N__16994),
            .I(N__16977));
    LocalMux I__3653 (
            .O(N__16989),
            .I(N__16974));
    Span4Mux_h I__3652 (
            .O(N__16986),
            .I(N__16971));
    InMux I__3651 (
            .O(N__16985),
            .I(N__16968));
    LocalMux I__3650 (
            .O(N__16982),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__3649 (
            .O(N__16977),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv12 I__3648 (
            .O(N__16974),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__3647 (
            .O(N__16971),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__3646 (
            .O(N__16968),
            .I(\Lab_UT.di_Mones_0 ));
    InMux I__3645 (
            .O(N__16957),
            .I(N__16950));
    InMux I__3644 (
            .O(N__16956),
            .I(N__16945));
    InMux I__3643 (
            .O(N__16955),
            .I(N__16945));
    InMux I__3642 (
            .O(N__16954),
            .I(N__16942));
    CascadeMux I__3641 (
            .O(N__16953),
            .I(N__16938));
    LocalMux I__3640 (
            .O(N__16950),
            .I(N__16931));
    LocalMux I__3639 (
            .O(N__16945),
            .I(N__16931));
    LocalMux I__3638 (
            .O(N__16942),
            .I(N__16931));
    InMux I__3637 (
            .O(N__16941),
            .I(N__16928));
    InMux I__3636 (
            .O(N__16938),
            .I(N__16925));
    Span4Mux_v I__3635 (
            .O(N__16931),
            .I(N__16922));
    LocalMux I__3634 (
            .O(N__16928),
            .I(N__16919));
    LocalMux I__3633 (
            .O(N__16925),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3632 (
            .O(N__16922),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3631 (
            .O(N__16919),
            .I(\Lab_UT.LdMones ));
    InMux I__3630 (
            .O(N__16912),
            .I(N__16901));
    InMux I__3629 (
            .O(N__16911),
            .I(N__16901));
    InMux I__3628 (
            .O(N__16910),
            .I(N__16890));
    InMux I__3627 (
            .O(N__16909),
            .I(N__16890));
    InMux I__3626 (
            .O(N__16908),
            .I(N__16890));
    InMux I__3625 (
            .O(N__16907),
            .I(N__16890));
    InMux I__3624 (
            .O(N__16906),
            .I(N__16890));
    LocalMux I__3623 (
            .O(N__16901),
            .I(\Lab_UT.sec2_0 ));
    LocalMux I__3622 (
            .O(N__16890),
            .I(\Lab_UT.sec2_0 ));
    CascadeMux I__3621 (
            .O(N__16885),
            .I(N__16878));
    CascadeMux I__3620 (
            .O(N__16884),
            .I(N__16875));
    CascadeMux I__3619 (
            .O(N__16883),
            .I(N__16871));
    CascadeMux I__3618 (
            .O(N__16882),
            .I(N__16867));
    InMux I__3617 (
            .O(N__16881),
            .I(N__16862));
    InMux I__3616 (
            .O(N__16878),
            .I(N__16862));
    InMux I__3615 (
            .O(N__16875),
            .I(N__16851));
    InMux I__3614 (
            .O(N__16874),
            .I(N__16851));
    InMux I__3613 (
            .O(N__16871),
            .I(N__16851));
    InMux I__3612 (
            .O(N__16870),
            .I(N__16851));
    InMux I__3611 (
            .O(N__16867),
            .I(N__16851));
    LocalMux I__3610 (
            .O(N__16862),
            .I(\Lab_UT.sec2_3 ));
    LocalMux I__3609 (
            .O(N__16851),
            .I(\Lab_UT.sec2_3 ));
    CascadeMux I__3608 (
            .O(N__16846),
            .I(N__16841));
    CascadeMux I__3607 (
            .O(N__16845),
            .I(N__16837));
    InMux I__3606 (
            .O(N__16844),
            .I(N__16823));
    InMux I__3605 (
            .O(N__16841),
            .I(N__16823));
    InMux I__3604 (
            .O(N__16840),
            .I(N__16823));
    InMux I__3603 (
            .O(N__16837),
            .I(N__16823));
    InMux I__3602 (
            .O(N__16836),
            .I(N__16823));
    InMux I__3601 (
            .O(N__16835),
            .I(N__16818));
    InMux I__3600 (
            .O(N__16834),
            .I(N__16818));
    LocalMux I__3599 (
            .O(N__16823),
            .I(N__16815));
    LocalMux I__3598 (
            .O(N__16818),
            .I(\Lab_UT.sec2_1 ));
    Odrv4 I__3597 (
            .O(N__16815),
            .I(\Lab_UT.sec2_1 ));
    CascadeMux I__3596 (
            .O(N__16810),
            .I(N__16807));
    InMux I__3595 (
            .O(N__16807),
            .I(N__16796));
    InMux I__3594 (
            .O(N__16806),
            .I(N__16796));
    InMux I__3593 (
            .O(N__16805),
            .I(N__16785));
    InMux I__3592 (
            .O(N__16804),
            .I(N__16785));
    InMux I__3591 (
            .O(N__16803),
            .I(N__16785));
    InMux I__3590 (
            .O(N__16802),
            .I(N__16785));
    InMux I__3589 (
            .O(N__16801),
            .I(N__16785));
    LocalMux I__3588 (
            .O(N__16796),
            .I(\Lab_UT.sec2_2 ));
    LocalMux I__3587 (
            .O(N__16785),
            .I(\Lab_UT.sec2_2 ));
    InMux I__3586 (
            .O(N__16780),
            .I(N__16776));
    InMux I__3585 (
            .O(N__16779),
            .I(N__16773));
    LocalMux I__3584 (
            .O(N__16776),
            .I(N__16770));
    LocalMux I__3583 (
            .O(N__16773),
            .I(\uu2.bitmapZ0Z_314 ));
    Odrv12 I__3582 (
            .O(N__16770),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__3581 (
            .O(N__16765),
            .I(N__16762));
    LocalMux I__3580 (
            .O(N__16762),
            .I(N__16756));
    InMux I__3579 (
            .O(N__16761),
            .I(N__16753));
    InMux I__3578 (
            .O(N__16760),
            .I(N__16750));
    InMux I__3577 (
            .O(N__16759),
            .I(N__16747));
    Span4Mux_h I__3576 (
            .O(N__16756),
            .I(N__16744));
    LocalMux I__3575 (
            .O(N__16753),
            .I(N__16739));
    LocalMux I__3574 (
            .O(N__16750),
            .I(N__16739));
    LocalMux I__3573 (
            .O(N__16747),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__3572 (
            .O(N__16744),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv12 I__3571 (
            .O(N__16739),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    InMux I__3570 (
            .O(N__16732),
            .I(N__16726));
    InMux I__3569 (
            .O(N__16731),
            .I(N__16726));
    LocalMux I__3568 (
            .O(N__16726),
            .I(N__16723));
    Span4Mux_h I__3567 (
            .O(N__16723),
            .I(N__16720));
    Odrv4 I__3566 (
            .O(N__16720),
            .I(\uu2.bitmap_RNIM5E21Z0Z_314 ));
    InMux I__3565 (
            .O(N__16717),
            .I(N__16710));
    InMux I__3564 (
            .O(N__16716),
            .I(N__16703));
    InMux I__3563 (
            .O(N__16715),
            .I(N__16703));
    InMux I__3562 (
            .O(N__16714),
            .I(N__16703));
    InMux I__3561 (
            .O(N__16713),
            .I(N__16700));
    LocalMux I__3560 (
            .O(N__16710),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3559 (
            .O(N__16703),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3558 (
            .O(N__16700),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    InMux I__3557 (
            .O(N__16693),
            .I(N__16690));
    LocalMux I__3556 (
            .O(N__16690),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__3555 (
            .O(N__16687),
            .I(N__16684));
    LocalMux I__3554 (
            .O(N__16684),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__3553 (
            .O(N__16681),
            .I(N__16678));
    LocalMux I__3552 (
            .O(N__16678),
            .I(\uu2.N_152 ));
    InMux I__3551 (
            .O(N__16675),
            .I(N__16672));
    LocalMux I__3550 (
            .O(N__16672),
            .I(N__16668));
    InMux I__3549 (
            .O(N__16671),
            .I(N__16665));
    Span4Mux_h I__3548 (
            .O(N__16668),
            .I(N__16662));
    LocalMux I__3547 (
            .O(N__16665),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    Odrv4 I__3546 (
            .O(N__16662),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__3545 (
            .O(N__16657),
            .I(N__16651));
    InMux I__3544 (
            .O(N__16656),
            .I(N__16651));
    LocalMux I__3543 (
            .O(N__16651),
            .I(N__16647));
    InMux I__3542 (
            .O(N__16650),
            .I(N__16644));
    Span4Mux_v I__3541 (
            .O(N__16647),
            .I(N__16639));
    LocalMux I__3540 (
            .O(N__16644),
            .I(N__16639));
    Odrv4 I__3539 (
            .O(N__16639),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    InMux I__3538 (
            .O(N__16636),
            .I(N__16628));
    InMux I__3537 (
            .O(N__16635),
            .I(N__16625));
    CascadeMux I__3536 (
            .O(N__16634),
            .I(N__16621));
    InMux I__3535 (
            .O(N__16633),
            .I(N__16614));
    InMux I__3534 (
            .O(N__16632),
            .I(N__16614));
    InMux I__3533 (
            .O(N__16631),
            .I(N__16614));
    LocalMux I__3532 (
            .O(N__16628),
            .I(N__16611));
    LocalMux I__3531 (
            .O(N__16625),
            .I(N__16608));
    InMux I__3530 (
            .O(N__16624),
            .I(N__16605));
    InMux I__3529 (
            .O(N__16621),
            .I(N__16602));
    LocalMux I__3528 (
            .O(N__16614),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__3527 (
            .O(N__16611),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__3526 (
            .O(N__16608),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__3525 (
            .O(N__16605),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__3524 (
            .O(N__16602),
            .I(\Lab_UT.di_Mtens_1 ));
    InMux I__3523 (
            .O(N__16591),
            .I(N__16587));
    InMux I__3522 (
            .O(N__16590),
            .I(N__16583));
    LocalMux I__3521 (
            .O(N__16587),
            .I(N__16580));
    InMux I__3520 (
            .O(N__16586),
            .I(N__16577));
    LocalMux I__3519 (
            .O(N__16583),
            .I(N__16574));
    Span4Mux_v I__3518 (
            .O(N__16580),
            .I(N__16569));
    LocalMux I__3517 (
            .O(N__16577),
            .I(N__16569));
    Odrv4 I__3516 (
            .O(N__16574),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv4 I__3515 (
            .O(N__16569),
            .I(\Lab_UT.di_AMtens_1 ));
    InMux I__3514 (
            .O(N__16564),
            .I(N__16561));
    LocalMux I__3513 (
            .O(N__16561),
            .I(N__16552));
    InMux I__3512 (
            .O(N__16560),
            .I(N__16539));
    InMux I__3511 (
            .O(N__16559),
            .I(N__16539));
    InMux I__3510 (
            .O(N__16558),
            .I(N__16539));
    InMux I__3509 (
            .O(N__16557),
            .I(N__16539));
    InMux I__3508 (
            .O(N__16556),
            .I(N__16539));
    InMux I__3507 (
            .O(N__16555),
            .I(N__16539));
    Span4Mux_h I__3506 (
            .O(N__16552),
            .I(N__16536));
    LocalMux I__3505 (
            .O(N__16539),
            .I(N__16533));
    Odrv4 I__3504 (
            .O(N__16536),
            .I(\Lab_UT.min1_1 ));
    Odrv4 I__3503 (
            .O(N__16533),
            .I(\Lab_UT.min1_1 ));
    CascadeMux I__3502 (
            .O(N__16528),
            .I(N__16525));
    InMux I__3501 (
            .O(N__16525),
            .I(N__16522));
    LocalMux I__3500 (
            .O(N__16522),
            .I(\Lab_UT.didp.countrce4.un13_qPone ));
    InMux I__3499 (
            .O(N__16519),
            .I(N__16516));
    LocalMux I__3498 (
            .O(N__16516),
            .I(\Lab_UT.didp.countrce4.q_5_2 ));
    InMux I__3497 (
            .O(N__16513),
            .I(N__16510));
    LocalMux I__3496 (
            .O(N__16510),
            .I(N__16507));
    Span4Mux_h I__3495 (
            .O(N__16507),
            .I(N__16504));
    Odrv4 I__3494 (
            .O(N__16504),
            .I(\uu2.bitmap_pmux_20_ns_1 ));
    InMux I__3493 (
            .O(N__16501),
            .I(N__16498));
    LocalMux I__3492 (
            .O(N__16498),
            .I(N__16495));
    Odrv4 I__3491 (
            .O(N__16495),
            .I(\uu2.bitmapZ0Z_162 ));
    InMux I__3490 (
            .O(N__16492),
            .I(N__16489));
    LocalMux I__3489 (
            .O(N__16489),
            .I(\uu2.bitmapZ0Z_290 ));
    InMux I__3488 (
            .O(N__16486),
            .I(N__16483));
    LocalMux I__3487 (
            .O(N__16483),
            .I(\uu2.bitmapZ0Z_34 ));
    CascadeMux I__3486 (
            .O(N__16480),
            .I(N__16477));
    InMux I__3485 (
            .O(N__16477),
            .I(N__16474));
    LocalMux I__3484 (
            .O(N__16474),
            .I(N__16471));
    Odrv4 I__3483 (
            .O(N__16471),
            .I(\uu2.bitmap_pmux_26_bm_1 ));
    CascadeMux I__3482 (
            .O(N__16468),
            .I(N__16464));
    CascadeMux I__3481 (
            .O(N__16467),
            .I(N__16459));
    InMux I__3480 (
            .O(N__16464),
            .I(N__16454));
    InMux I__3479 (
            .O(N__16463),
            .I(N__16451));
    InMux I__3478 (
            .O(N__16462),
            .I(N__16446));
    InMux I__3477 (
            .O(N__16459),
            .I(N__16446));
    InMux I__3476 (
            .O(N__16458),
            .I(N__16441));
    InMux I__3475 (
            .O(N__16457),
            .I(N__16441));
    LocalMux I__3474 (
            .O(N__16454),
            .I(N__16436));
    LocalMux I__3473 (
            .O(N__16451),
            .I(N__16436));
    LocalMux I__3472 (
            .O(N__16446),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3471 (
            .O(N__16441),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv12 I__3470 (
            .O(N__16436),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__3469 (
            .O(N__16429),
            .I(N__16426));
    LocalMux I__3468 (
            .O(N__16426),
            .I(N__16423));
    Odrv4 I__3467 (
            .O(N__16423),
            .I(\uu2.bitmap_RNIP2JO1Z0Z_34 ));
    InMux I__3466 (
            .O(N__16420),
            .I(N__16411));
    InMux I__3465 (
            .O(N__16419),
            .I(N__16398));
    InMux I__3464 (
            .O(N__16418),
            .I(N__16398));
    InMux I__3463 (
            .O(N__16417),
            .I(N__16398));
    InMux I__3462 (
            .O(N__16416),
            .I(N__16398));
    InMux I__3461 (
            .O(N__16415),
            .I(N__16398));
    InMux I__3460 (
            .O(N__16414),
            .I(N__16398));
    LocalMux I__3459 (
            .O(N__16411),
            .I(N__16395));
    LocalMux I__3458 (
            .O(N__16398),
            .I(\Lab_UT.min1_0 ));
    Odrv4 I__3457 (
            .O(N__16395),
            .I(\Lab_UT.min1_0 ));
    CascadeMux I__3456 (
            .O(N__16390),
            .I(N__16384));
    CascadeMux I__3455 (
            .O(N__16389),
            .I(N__16380));
    CascadeMux I__3454 (
            .O(N__16388),
            .I(N__16376));
    CascadeMux I__3453 (
            .O(N__16387),
            .I(N__16372));
    InMux I__3452 (
            .O(N__16384),
            .I(N__16359));
    InMux I__3451 (
            .O(N__16383),
            .I(N__16359));
    InMux I__3450 (
            .O(N__16380),
            .I(N__16359));
    InMux I__3449 (
            .O(N__16379),
            .I(N__16359));
    InMux I__3448 (
            .O(N__16376),
            .I(N__16359));
    InMux I__3447 (
            .O(N__16375),
            .I(N__16359));
    InMux I__3446 (
            .O(N__16372),
            .I(N__16356));
    LocalMux I__3445 (
            .O(N__16359),
            .I(N__16353));
    LocalMux I__3444 (
            .O(N__16356),
            .I(N__16350));
    Odrv4 I__3443 (
            .O(N__16353),
            .I(\Lab_UT.min1_3 ));
    Odrv12 I__3442 (
            .O(N__16350),
            .I(\Lab_UT.min1_3 ));
    InMux I__3441 (
            .O(N__16345),
            .I(N__16342));
    LocalMux I__3440 (
            .O(N__16342),
            .I(N__16339));
    Span4Mux_h I__3439 (
            .O(N__16339),
            .I(N__16336));
    Odrv4 I__3438 (
            .O(N__16336),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__3437 (
            .O(N__16333),
            .I(N__16326));
    InMux I__3436 (
            .O(N__16332),
            .I(N__16326));
    InMux I__3435 (
            .O(N__16331),
            .I(N__16318));
    LocalMux I__3434 (
            .O(N__16326),
            .I(N__16315));
    CascadeMux I__3433 (
            .O(N__16325),
            .I(N__16312));
    InMux I__3432 (
            .O(N__16324),
            .I(N__16306));
    InMux I__3431 (
            .O(N__16323),
            .I(N__16299));
    InMux I__3430 (
            .O(N__16322),
            .I(N__16299));
    InMux I__3429 (
            .O(N__16321),
            .I(N__16299));
    LocalMux I__3428 (
            .O(N__16318),
            .I(N__16294));
    Span4Mux_v I__3427 (
            .O(N__16315),
            .I(N__16294));
    InMux I__3426 (
            .O(N__16312),
            .I(N__16289));
    InMux I__3425 (
            .O(N__16311),
            .I(N__16289));
    InMux I__3424 (
            .O(N__16310),
            .I(N__16286));
    InMux I__3423 (
            .O(N__16309),
            .I(N__16283));
    LocalMux I__3422 (
            .O(N__16306),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3421 (
            .O(N__16299),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3420 (
            .O(N__16294),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3419 (
            .O(N__16289),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3418 (
            .O(N__16286),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3417 (
            .O(N__16283),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__3416 (
            .O(N__16270),
            .I(N__16267));
    LocalMux I__3415 (
            .O(N__16267),
            .I(\uu2.bitmapZ0Z_218 ));
    CascadeMux I__3414 (
            .O(N__16264),
            .I(N__16259));
    CascadeMux I__3413 (
            .O(N__16263),
            .I(N__16256));
    CascadeMux I__3412 (
            .O(N__16262),
            .I(N__16252));
    InMux I__3411 (
            .O(N__16259),
            .I(N__16246));
    InMux I__3410 (
            .O(N__16256),
            .I(N__16237));
    InMux I__3409 (
            .O(N__16255),
            .I(N__16237));
    InMux I__3408 (
            .O(N__16252),
            .I(N__16237));
    InMux I__3407 (
            .O(N__16251),
            .I(N__16237));
    CascadeMux I__3406 (
            .O(N__16250),
            .I(N__16231));
    InMux I__3405 (
            .O(N__16249),
            .I(N__16228));
    LocalMux I__3404 (
            .O(N__16246),
            .I(N__16223));
    LocalMux I__3403 (
            .O(N__16237),
            .I(N__16223));
    InMux I__3402 (
            .O(N__16236),
            .I(N__16216));
    InMux I__3401 (
            .O(N__16235),
            .I(N__16216));
    InMux I__3400 (
            .O(N__16234),
            .I(N__16216));
    InMux I__3399 (
            .O(N__16231),
            .I(N__16213));
    LocalMux I__3398 (
            .O(N__16228),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3397 (
            .O(N__16223),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3396 (
            .O(N__16216),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3395 (
            .O(N__16213),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__3394 (
            .O(N__16204),
            .I(N__16201));
    LocalMux I__3393 (
            .O(N__16201),
            .I(\uu2.bitmapZ0Z_90 ));
    InMux I__3392 (
            .O(N__16198),
            .I(N__16195));
    LocalMux I__3391 (
            .O(N__16195),
            .I(N__16192));
    Odrv4 I__3390 (
            .O(N__16192),
            .I(\uu2.bitmap_pmux_19_ns_1 ));
    InMux I__3389 (
            .O(N__16189),
            .I(N__16182));
    InMux I__3388 (
            .O(N__16188),
            .I(N__16177));
    InMux I__3387 (
            .O(N__16187),
            .I(N__16177));
    InMux I__3386 (
            .O(N__16186),
            .I(N__16172));
    InMux I__3385 (
            .O(N__16185),
            .I(N__16172));
    LocalMux I__3384 (
            .O(N__16182),
            .I(N__16167));
    LocalMux I__3383 (
            .O(N__16177),
            .I(N__16167));
    LocalMux I__3382 (
            .O(N__16172),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__3381 (
            .O(N__16167),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__3380 (
            .O(N__16162),
            .I(\uu2.un3_w_addr_user_4_cascade_ ));
    InMux I__3379 (
            .O(N__16159),
            .I(N__16156));
    LocalMux I__3378 (
            .O(N__16156),
            .I(\uu2.un3_w_addr_user_5 ));
    InMux I__3377 (
            .O(N__16153),
            .I(N__16147));
    InMux I__3376 (
            .O(N__16152),
            .I(N__16147));
    LocalMux I__3375 (
            .O(N__16147),
            .I(N__16144));
    Span4Mux_h I__3374 (
            .O(N__16144),
            .I(N__16141));
    Odrv4 I__3373 (
            .O(N__16141),
            .I(\uu2.un3_w_addr_user ));
    InMux I__3372 (
            .O(N__16138),
            .I(N__16132));
    InMux I__3371 (
            .O(N__16137),
            .I(N__16129));
    CascadeMux I__3370 (
            .O(N__16136),
            .I(N__16123));
    CascadeMux I__3369 (
            .O(N__16135),
            .I(N__16120));
    LocalMux I__3368 (
            .O(N__16132),
            .I(N__16116));
    LocalMux I__3367 (
            .O(N__16129),
            .I(N__16113));
    CascadeMux I__3366 (
            .O(N__16128),
            .I(N__16108));
    InMux I__3365 (
            .O(N__16127),
            .I(N__16103));
    InMux I__3364 (
            .O(N__16126),
            .I(N__16103));
    InMux I__3363 (
            .O(N__16123),
            .I(N__16098));
    InMux I__3362 (
            .O(N__16120),
            .I(N__16098));
    InMux I__3361 (
            .O(N__16119),
            .I(N__16095));
    Span4Mux_v I__3360 (
            .O(N__16116),
            .I(N__16092));
    Span4Mux_s1_v I__3359 (
            .O(N__16113),
            .I(N__16089));
    InMux I__3358 (
            .O(N__16112),
            .I(N__16084));
    InMux I__3357 (
            .O(N__16111),
            .I(N__16084));
    InMux I__3356 (
            .O(N__16108),
            .I(N__16081));
    LocalMux I__3355 (
            .O(N__16103),
            .I(N__16072));
    LocalMux I__3354 (
            .O(N__16098),
            .I(N__16072));
    LocalMux I__3353 (
            .O(N__16095),
            .I(N__16072));
    Span4Mux_s1_v I__3352 (
            .O(N__16092),
            .I(N__16072));
    Odrv4 I__3351 (
            .O(N__16089),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3350 (
            .O(N__16084),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3349 (
            .O(N__16081),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__3348 (
            .O(N__16072),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    CascadeMux I__3347 (
            .O(N__16063),
            .I(N__16060));
    InMux I__3346 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__3345 (
            .O(N__16057),
            .I(N__16054));
    Odrv12 I__3344 (
            .O(N__16054),
            .I(\uu2.mem0.w_addr_3 ));
    InMux I__3343 (
            .O(N__16051),
            .I(N__16044));
    InMux I__3342 (
            .O(N__16050),
            .I(N__16041));
    InMux I__3341 (
            .O(N__16049),
            .I(N__16036));
    InMux I__3340 (
            .O(N__16048),
            .I(N__16036));
    InMux I__3339 (
            .O(N__16047),
            .I(N__16033));
    LocalMux I__3338 (
            .O(N__16044),
            .I(N__16026));
    LocalMux I__3337 (
            .O(N__16041),
            .I(N__16026));
    LocalMux I__3336 (
            .O(N__16036),
            .I(N__16026));
    LocalMux I__3335 (
            .O(N__16033),
            .I(N__16023));
    Odrv12 I__3334 (
            .O(N__16026),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__3333 (
            .O(N__16023),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__3332 (
            .O(N__16018),
            .I(N__16015));
    InMux I__3331 (
            .O(N__16015),
            .I(N__16009));
    InMux I__3330 (
            .O(N__16014),
            .I(N__16004));
    InMux I__3329 (
            .O(N__16013),
            .I(N__16004));
    InMux I__3328 (
            .O(N__16012),
            .I(N__16001));
    LocalMux I__3327 (
            .O(N__16009),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__3326 (
            .O(N__16004),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__3325 (
            .O(N__16001),
            .I(\uu2.w_addr_userZ0Z_7 ));
    CascadeMux I__3324 (
            .O(N__15994),
            .I(N__15990));
    InMux I__3323 (
            .O(N__15993),
            .I(N__15979));
    InMux I__3322 (
            .O(N__15990),
            .I(N__15979));
    InMux I__3321 (
            .O(N__15989),
            .I(N__15979));
    InMux I__3320 (
            .O(N__15988),
            .I(N__15979));
    LocalMux I__3319 (
            .O(N__15979),
            .I(\uu2.w_addr_userZ0Z_3 ));
    InMux I__3318 (
            .O(N__15976),
            .I(N__15973));
    LocalMux I__3317 (
            .O(N__15973),
            .I(N__15970));
    Span4Mux_v I__3316 (
            .O(N__15970),
            .I(N__15963));
    InMux I__3315 (
            .O(N__15969),
            .I(N__15954));
    InMux I__3314 (
            .O(N__15968),
            .I(N__15954));
    InMux I__3313 (
            .O(N__15967),
            .I(N__15954));
    InMux I__3312 (
            .O(N__15966),
            .I(N__15951));
    Span4Mux_h I__3311 (
            .O(N__15963),
            .I(N__15948));
    InMux I__3310 (
            .O(N__15962),
            .I(N__15943));
    InMux I__3309 (
            .O(N__15961),
            .I(N__15943));
    LocalMux I__3308 (
            .O(N__15954),
            .I(N__15940));
    LocalMux I__3307 (
            .O(N__15951),
            .I(N__15935));
    Span4Mux_v I__3306 (
            .O(N__15948),
            .I(N__15935));
    LocalMux I__3305 (
            .O(N__15943),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__3304 (
            .O(N__15940),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__3303 (
            .O(N__15935),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__3302 (
            .O(N__15928),
            .I(N__15924));
    InMux I__3301 (
            .O(N__15927),
            .I(N__15916));
    InMux I__3300 (
            .O(N__15924),
            .I(N__15916));
    InMux I__3299 (
            .O(N__15923),
            .I(N__15916));
    LocalMux I__3298 (
            .O(N__15916),
            .I(N__15912));
    InMux I__3297 (
            .O(N__15915),
            .I(N__15909));
    Odrv4 I__3296 (
            .O(N__15912),
            .I(\uu2.un404_ci ));
    LocalMux I__3295 (
            .O(N__15909),
            .I(\uu2.un404_ci ));
    CascadeMux I__3294 (
            .O(N__15904),
            .I(N__15899));
    InMux I__3293 (
            .O(N__15903),
            .I(N__15894));
    InMux I__3292 (
            .O(N__15902),
            .I(N__15894));
    InMux I__3291 (
            .O(N__15899),
            .I(N__15891));
    LocalMux I__3290 (
            .O(N__15894),
            .I(N__15888));
    LocalMux I__3289 (
            .O(N__15891),
            .I(N__15885));
    Odrv4 I__3288 (
            .O(N__15888),
            .I(\uu2.un426_ci_3 ));
    Odrv4 I__3287 (
            .O(N__15885),
            .I(\uu2.un426_ci_3 ));
    CascadeMux I__3286 (
            .O(N__15880),
            .I(\uu2.un404_ci_cascade_ ));
    InMux I__3285 (
            .O(N__15877),
            .I(N__15874));
    LocalMux I__3284 (
            .O(N__15874),
            .I(\uu2.vbuf_w_addr_user.un448_ci_0 ));
    InMux I__3283 (
            .O(N__15871),
            .I(N__15868));
    LocalMux I__3282 (
            .O(N__15868),
            .I(N__15863));
    InMux I__3281 (
            .O(N__15867),
            .I(N__15858));
    InMux I__3280 (
            .O(N__15866),
            .I(N__15858));
    Odrv12 I__3279 (
            .O(N__15863),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__3278 (
            .O(N__15858),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CEMux I__3277 (
            .O(N__15853),
            .I(N__15850));
    LocalMux I__3276 (
            .O(N__15850),
            .I(N__15847));
    Sp12to4 I__3275 (
            .O(N__15847),
            .I(N__15844));
    Odrv12 I__3274 (
            .O(N__15844),
            .I(\uu2.un28_w_addr_user_i_0 ));
    SRMux I__3273 (
            .O(N__15841),
            .I(N__15838));
    LocalMux I__3272 (
            .O(N__15838),
            .I(N__15835));
    Span4Mux_s0_v I__3271 (
            .O(N__15835),
            .I(N__15831));
    SRMux I__3270 (
            .O(N__15834),
            .I(N__15828));
    Span4Mux_h I__3269 (
            .O(N__15831),
            .I(N__15823));
    LocalMux I__3268 (
            .O(N__15828),
            .I(N__15823));
    Span4Mux_s0_v I__3267 (
            .O(N__15823),
            .I(N__15819));
    InMux I__3266 (
            .O(N__15822),
            .I(N__15816));
    Odrv4 I__3265 (
            .O(N__15819),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_4 ));
    LocalMux I__3264 (
            .O(N__15816),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_4 ));
    InMux I__3263 (
            .O(N__15811),
            .I(N__15808));
    LocalMux I__3262 (
            .O(N__15808),
            .I(\uu2.bitmapZ0Z_194 ));
    InMux I__3261 (
            .O(N__15805),
            .I(N__15802));
    LocalMux I__3260 (
            .O(N__15802),
            .I(\uu2.bitmapZ0Z_66 ));
    CascadeMux I__3259 (
            .O(N__15799),
            .I(N__15796));
    InMux I__3258 (
            .O(N__15796),
            .I(N__15790));
    InMux I__3257 (
            .O(N__15795),
            .I(N__15790));
    LocalMux I__3256 (
            .O(N__15790),
            .I(N__15780));
    InMux I__3255 (
            .O(N__15789),
            .I(N__15775));
    InMux I__3254 (
            .O(N__15788),
            .I(N__15775));
    CascadeMux I__3253 (
            .O(N__15787),
            .I(N__15772));
    InMux I__3252 (
            .O(N__15786),
            .I(N__15769));
    CascadeMux I__3251 (
            .O(N__15785),
            .I(N__15766));
    CascadeMux I__3250 (
            .O(N__15784),
            .I(N__15762));
    InMux I__3249 (
            .O(N__15783),
            .I(N__15759));
    Span4Mux_v I__3248 (
            .O(N__15780),
            .I(N__15754));
    LocalMux I__3247 (
            .O(N__15775),
            .I(N__15754));
    InMux I__3246 (
            .O(N__15772),
            .I(N__15751));
    LocalMux I__3245 (
            .O(N__15769),
            .I(N__15748));
    InMux I__3244 (
            .O(N__15766),
            .I(N__15745));
    InMux I__3243 (
            .O(N__15765),
            .I(N__15740));
    InMux I__3242 (
            .O(N__15762),
            .I(N__15740));
    LocalMux I__3241 (
            .O(N__15759),
            .I(N__15737));
    Span4Mux_h I__3240 (
            .O(N__15754),
            .I(N__15734));
    LocalMux I__3239 (
            .O(N__15751),
            .I(N__15727));
    Span4Mux_h I__3238 (
            .O(N__15748),
            .I(N__15727));
    LocalMux I__3237 (
            .O(N__15745),
            .I(N__15727));
    LocalMux I__3236 (
            .O(N__15740),
            .I(N__15724));
    Odrv12 I__3235 (
            .O(N__15737),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__3234 (
            .O(N__15734),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__3233 (
            .O(N__15727),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__3232 (
            .O(N__15724),
            .I(bu_rx_data_2_rep1));
    CascadeMux I__3231 (
            .O(N__15715),
            .I(N__15712));
    InMux I__3230 (
            .O(N__15712),
            .I(N__15705));
    InMux I__3229 (
            .O(N__15711),
            .I(N__15700));
    InMux I__3228 (
            .O(N__15710),
            .I(N__15700));
    InMux I__3227 (
            .O(N__15709),
            .I(N__15695));
    InMux I__3226 (
            .O(N__15708),
            .I(N__15692));
    LocalMux I__3225 (
            .O(N__15705),
            .I(N__15687));
    LocalMux I__3224 (
            .O(N__15700),
            .I(N__15687));
    InMux I__3223 (
            .O(N__15699),
            .I(N__15682));
    InMux I__3222 (
            .O(N__15698),
            .I(N__15682));
    LocalMux I__3221 (
            .O(N__15695),
            .I(N__15679));
    LocalMux I__3220 (
            .O(N__15692),
            .I(N__15676));
    Span4Mux_h I__3219 (
            .O(N__15687),
            .I(N__15673));
    LocalMux I__3218 (
            .O(N__15682),
            .I(N__15670));
    Odrv4 I__3217 (
            .O(N__15679),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__3216 (
            .O(N__15676),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__3215 (
            .O(N__15673),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__3214 (
            .O(N__15670),
            .I(bu_rx_data_0_rep1));
    CascadeMux I__3213 (
            .O(N__15661),
            .I(N__15658));
    InMux I__3212 (
            .O(N__15658),
            .I(N__15655));
    LocalMux I__3211 (
            .O(N__15655),
            .I(N__15652));
    Odrv4 I__3210 (
            .O(N__15652),
            .I(G_6_0_a6_3_3));
    InMux I__3209 (
            .O(N__15649),
            .I(N__15642));
    InMux I__3208 (
            .O(N__15648),
            .I(N__15637));
    InMux I__3207 (
            .O(N__15647),
            .I(N__15637));
    InMux I__3206 (
            .O(N__15646),
            .I(N__15632));
    InMux I__3205 (
            .O(N__15645),
            .I(N__15632));
    LocalMux I__3204 (
            .O(N__15642),
            .I(buart__rx_shifter_fast_4));
    LocalMux I__3203 (
            .O(N__15637),
            .I(buart__rx_shifter_fast_4));
    LocalMux I__3202 (
            .O(N__15632),
            .I(buart__rx_shifter_fast_4));
    CascadeMux I__3201 (
            .O(N__15625),
            .I(N__15618));
    InMux I__3200 (
            .O(N__15624),
            .I(N__15615));
    InMux I__3199 (
            .O(N__15623),
            .I(N__15606));
    InMux I__3198 (
            .O(N__15622),
            .I(N__15606));
    InMux I__3197 (
            .O(N__15621),
            .I(N__15606));
    InMux I__3196 (
            .O(N__15618),
            .I(N__15606));
    LocalMux I__3195 (
            .O(N__15615),
            .I(bu_rx_data_7_rep1));
    LocalMux I__3194 (
            .O(N__15606),
            .I(bu_rx_data_7_rep1));
    InMux I__3193 (
            .O(N__15601),
            .I(N__15594));
    InMux I__3192 (
            .O(N__15600),
            .I(N__15594));
    InMux I__3191 (
            .O(N__15599),
            .I(N__15591));
    LocalMux I__3190 (
            .O(N__15594),
            .I(N__15586));
    LocalMux I__3189 (
            .O(N__15591),
            .I(N__15586));
    Span4Mux_v I__3188 (
            .O(N__15586),
            .I(N__15582));
    InMux I__3187 (
            .O(N__15585),
            .I(N__15579));
    Span4Mux_v I__3186 (
            .O(N__15582),
            .I(N__15576));
    LocalMux I__3185 (
            .O(N__15579),
            .I(N__15573));
    Span4Mux_v I__3184 (
            .O(N__15576),
            .I(N__15568));
    Span4Mux_s3_v I__3183 (
            .O(N__15573),
            .I(N__15568));
    Odrv4 I__3182 (
            .O(N__15568),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    CascadeMux I__3181 (
            .O(N__15565),
            .I(N__15555));
    InMux I__3180 (
            .O(N__15564),
            .I(N__15550));
    InMux I__3179 (
            .O(N__15563),
            .I(N__15547));
    InMux I__3178 (
            .O(N__15562),
            .I(N__15544));
    InMux I__3177 (
            .O(N__15561),
            .I(N__15541));
    InMux I__3176 (
            .O(N__15560),
            .I(N__15536));
    InMux I__3175 (
            .O(N__15559),
            .I(N__15536));
    InMux I__3174 (
            .O(N__15558),
            .I(N__15533));
    InMux I__3173 (
            .O(N__15555),
            .I(N__15526));
    InMux I__3172 (
            .O(N__15554),
            .I(N__15526));
    InMux I__3171 (
            .O(N__15553),
            .I(N__15526));
    LocalMux I__3170 (
            .O(N__15550),
            .I(N__15521));
    LocalMux I__3169 (
            .O(N__15547),
            .I(N__15512));
    LocalMux I__3168 (
            .O(N__15544),
            .I(N__15512));
    LocalMux I__3167 (
            .O(N__15541),
            .I(N__15512));
    LocalMux I__3166 (
            .O(N__15536),
            .I(N__15512));
    LocalMux I__3165 (
            .O(N__15533),
            .I(N__15507));
    LocalMux I__3164 (
            .O(N__15526),
            .I(N__15507));
    InMux I__3163 (
            .O(N__15525),
            .I(N__15504));
    InMux I__3162 (
            .O(N__15524),
            .I(N__15501));
    Span4Mux_h I__3161 (
            .O(N__15521),
            .I(N__15498));
    Span4Mux_h I__3160 (
            .O(N__15512),
            .I(N__15495));
    Span4Mux_h I__3159 (
            .O(N__15507),
            .I(N__15492));
    LocalMux I__3158 (
            .O(N__15504),
            .I(bu_rx_data_7));
    LocalMux I__3157 (
            .O(N__15501),
            .I(bu_rx_data_7));
    Odrv4 I__3156 (
            .O(N__15498),
            .I(bu_rx_data_7));
    Odrv4 I__3155 (
            .O(N__15495),
            .I(bu_rx_data_7));
    Odrv4 I__3154 (
            .O(N__15492),
            .I(bu_rx_data_7));
    CEMux I__3153 (
            .O(N__15481),
            .I(N__15454));
    CEMux I__3152 (
            .O(N__15480),
            .I(N__15454));
    CEMux I__3151 (
            .O(N__15479),
            .I(N__15454));
    CEMux I__3150 (
            .O(N__15478),
            .I(N__15454));
    CEMux I__3149 (
            .O(N__15477),
            .I(N__15454));
    CEMux I__3148 (
            .O(N__15476),
            .I(N__15454));
    CEMux I__3147 (
            .O(N__15475),
            .I(N__15454));
    CEMux I__3146 (
            .O(N__15474),
            .I(N__15454));
    CEMux I__3145 (
            .O(N__15473),
            .I(N__15454));
    GlobalMux I__3144 (
            .O(N__15454),
            .I(N__15451));
    gio2CtrlBuf I__3143 (
            .O(N__15451),
            .I(\buart.Z_rx.sample_g ));
    CascadeMux I__3142 (
            .O(N__15448),
            .I(N__15445));
    InMux I__3141 (
            .O(N__15445),
            .I(N__15440));
    InMux I__3140 (
            .O(N__15444),
            .I(N__15434));
    InMux I__3139 (
            .O(N__15443),
            .I(N__15434));
    LocalMux I__3138 (
            .O(N__15440),
            .I(N__15431));
    InMux I__3137 (
            .O(N__15439),
            .I(N__15428));
    LocalMux I__3136 (
            .O(N__15434),
            .I(N__15425));
    Span4Mux_h I__3135 (
            .O(N__15431),
            .I(N__15422));
    LocalMux I__3134 (
            .O(N__15428),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__3133 (
            .O(N__15425),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__3132 (
            .O(N__15422),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__3131 (
            .O(N__15415),
            .I(\Lab_UT.dictrl.m22_xZ0Z1_cascade_ ));
    CascadeMux I__3130 (
            .O(N__15412),
            .I(\Lab_UT.dictrl.N_72_mux_cascade_ ));
    InMux I__3129 (
            .O(N__15409),
            .I(N__15406));
    LocalMux I__3128 (
            .O(N__15406),
            .I(N__15400));
    InMux I__3127 (
            .O(N__15405),
            .I(N__15397));
    InMux I__3126 (
            .O(N__15404),
            .I(N__15394));
    InMux I__3125 (
            .O(N__15403),
            .I(N__15391));
    Span4Mux_s3_v I__3124 (
            .O(N__15400),
            .I(N__15379));
    LocalMux I__3123 (
            .O(N__15397),
            .I(N__15379));
    LocalMux I__3122 (
            .O(N__15394),
            .I(N__15372));
    LocalMux I__3121 (
            .O(N__15391),
            .I(N__15372));
    InMux I__3120 (
            .O(N__15390),
            .I(N__15369));
    InMux I__3119 (
            .O(N__15389),
            .I(N__15366));
    InMux I__3118 (
            .O(N__15388),
            .I(N__15361));
    InMux I__3117 (
            .O(N__15387),
            .I(N__15361));
    InMux I__3116 (
            .O(N__15386),
            .I(N__15354));
    InMux I__3115 (
            .O(N__15385),
            .I(N__15354));
    InMux I__3114 (
            .O(N__15384),
            .I(N__15354));
    Span4Mux_h I__3113 (
            .O(N__15379),
            .I(N__15351));
    InMux I__3112 (
            .O(N__15378),
            .I(N__15346));
    InMux I__3111 (
            .O(N__15377),
            .I(N__15346));
    Odrv4 I__3110 (
            .O(N__15372),
            .I(bu_rx_data_4));
    LocalMux I__3109 (
            .O(N__15369),
            .I(bu_rx_data_4));
    LocalMux I__3108 (
            .O(N__15366),
            .I(bu_rx_data_4));
    LocalMux I__3107 (
            .O(N__15361),
            .I(bu_rx_data_4));
    LocalMux I__3106 (
            .O(N__15354),
            .I(bu_rx_data_4));
    Odrv4 I__3105 (
            .O(N__15351),
            .I(bu_rx_data_4));
    LocalMux I__3104 (
            .O(N__15346),
            .I(bu_rx_data_4));
    CascadeMux I__3103 (
            .O(N__15331),
            .I(N__15328));
    InMux I__3102 (
            .O(N__15328),
            .I(N__15324));
    CascadeMux I__3101 (
            .O(N__15327),
            .I(N__15321));
    LocalMux I__3100 (
            .O(N__15324),
            .I(N__15318));
    InMux I__3099 (
            .O(N__15321),
            .I(N__15315));
    Span4Mux_v I__3098 (
            .O(N__15318),
            .I(N__15312));
    LocalMux I__3097 (
            .O(N__15315),
            .I(bu_rx_data_fast_3));
    Odrv4 I__3096 (
            .O(N__15312),
            .I(bu_rx_data_fast_3));
    CascadeMux I__3095 (
            .O(N__15307),
            .I(N__15303));
    CascadeMux I__3094 (
            .O(N__15306),
            .I(N__15300));
    InMux I__3093 (
            .O(N__15303),
            .I(N__15294));
    InMux I__3092 (
            .O(N__15300),
            .I(N__15294));
    InMux I__3091 (
            .O(N__15299),
            .I(N__15291));
    LocalMux I__3090 (
            .O(N__15294),
            .I(N__15288));
    LocalMux I__3089 (
            .O(N__15291),
            .I(N__15285));
    Odrv4 I__3088 (
            .O(N__15288),
            .I(\Lab_UT.dictrl.m34Z0Z_1 ));
    Odrv4 I__3087 (
            .O(N__15285),
            .I(\Lab_UT.dictrl.m34Z0Z_1 ));
    CascadeMux I__3086 (
            .O(N__15280),
            .I(\Lab_UT.dictrl.g1_0_xZ0Z1_cascade_ ));
    InMux I__3085 (
            .O(N__15277),
            .I(N__15274));
    LocalMux I__3084 (
            .O(N__15274),
            .I(N__15271));
    Odrv4 I__3083 (
            .O(N__15271),
            .I(\Lab_UT.dictrl.g1_0_4 ));
    InMux I__3082 (
            .O(N__15268),
            .I(N__15265));
    LocalMux I__3081 (
            .O(N__15265),
            .I(\Lab_UT.dictrl.g0_5_3 ));
    CascadeMux I__3080 (
            .O(N__15262),
            .I(\Lab_UT.dictrl.g1_0_cascade_ ));
    InMux I__3079 (
            .O(N__15259),
            .I(N__15252));
    InMux I__3078 (
            .O(N__15258),
            .I(N__15252));
    CascadeMux I__3077 (
            .O(N__15257),
            .I(N__15249));
    LocalMux I__3076 (
            .O(N__15252),
            .I(N__15245));
    InMux I__3075 (
            .O(N__15249),
            .I(N__15242));
    InMux I__3074 (
            .O(N__15248),
            .I(N__15239));
    Odrv4 I__3073 (
            .O(N__15245),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    LocalMux I__3072 (
            .O(N__15242),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    LocalMux I__3071 (
            .O(N__15239),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    InMux I__3070 (
            .O(N__15232),
            .I(N__15229));
    LocalMux I__3069 (
            .O(N__15229),
            .I(\Lab_UT.dictrl.g0_5Z0Z_4 ));
    InMux I__3068 (
            .O(N__15226),
            .I(N__15220));
    InMux I__3067 (
            .O(N__15225),
            .I(N__15215));
    InMux I__3066 (
            .O(N__15224),
            .I(N__15215));
    InMux I__3065 (
            .O(N__15223),
            .I(N__15212));
    LocalMux I__3064 (
            .O(N__15220),
            .I(N__15207));
    LocalMux I__3063 (
            .O(N__15215),
            .I(N__15207));
    LocalMux I__3062 (
            .O(N__15212),
            .I(N__15202));
    Span4Mux_v I__3061 (
            .O(N__15207),
            .I(N__15202));
    Odrv4 I__3060 (
            .O(N__15202),
            .I(\Lab_UT.dictrl.next_state66_2 ));
    CascadeMux I__3059 (
            .O(N__15199),
            .I(N__15195));
    CascadeMux I__3058 (
            .O(N__15198),
            .I(N__15191));
    InMux I__3057 (
            .O(N__15195),
            .I(N__15188));
    InMux I__3056 (
            .O(N__15194),
            .I(N__15180));
    InMux I__3055 (
            .O(N__15191),
            .I(N__15177));
    LocalMux I__3054 (
            .O(N__15188),
            .I(N__15174));
    InMux I__3053 (
            .O(N__15187),
            .I(N__15169));
    InMux I__3052 (
            .O(N__15186),
            .I(N__15169));
    InMux I__3051 (
            .O(N__15185),
            .I(N__15162));
    InMux I__3050 (
            .O(N__15184),
            .I(N__15162));
    InMux I__3049 (
            .O(N__15183),
            .I(N__15162));
    LocalMux I__3048 (
            .O(N__15180),
            .I(N__15159));
    LocalMux I__3047 (
            .O(N__15177),
            .I(N__15152));
    Span4Mux_h I__3046 (
            .O(N__15174),
            .I(N__15152));
    LocalMux I__3045 (
            .O(N__15169),
            .I(N__15152));
    LocalMux I__3044 (
            .O(N__15162),
            .I(N__15149));
    Span4Mux_v I__3043 (
            .O(N__15159),
            .I(N__15146));
    Span4Mux_v I__3042 (
            .O(N__15152),
            .I(N__15143));
    Sp12to4 I__3041 (
            .O(N__15149),
            .I(N__15140));
    Odrv4 I__3040 (
            .O(N__15146),
            .I(\Lab_UT.dictrl.state_i_3_0 ));
    Odrv4 I__3039 (
            .O(N__15143),
            .I(\Lab_UT.dictrl.state_i_3_0 ));
    Odrv12 I__3038 (
            .O(N__15140),
            .I(\Lab_UT.dictrl.state_i_3_0 ));
    CascadeMux I__3037 (
            .O(N__15133),
            .I(N_5_cascade_));
    InMux I__3036 (
            .O(N__15130),
            .I(N__15127));
    LocalMux I__3035 (
            .O(N__15127),
            .I(N__15124));
    Span4Mux_h I__3034 (
            .O(N__15124),
            .I(N__15121));
    Odrv4 I__3033 (
            .O(N__15121),
            .I(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ));
    CascadeMux I__3032 (
            .O(N__15118),
            .I(\Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_ ));
    InMux I__3031 (
            .O(N__15115),
            .I(N__15111));
    InMux I__3030 (
            .O(N__15114),
            .I(N__15108));
    LocalMux I__3029 (
            .O(N__15111),
            .I(\Lab_UT.dictrl.N_67_mux ));
    LocalMux I__3028 (
            .O(N__15108),
            .I(\Lab_UT.dictrl.N_67_mux ));
    InMux I__3027 (
            .O(N__15103),
            .I(N__15100));
    LocalMux I__3026 (
            .O(N__15100),
            .I(N__15097));
    Odrv4 I__3025 (
            .O(N__15097),
            .I(\Lab_UT.dictrl.G_6_0_1_0 ));
    InMux I__3024 (
            .O(N__15094),
            .I(N__15091));
    LocalMux I__3023 (
            .O(N__15091),
            .I(\Lab_UT.dictrl.N_12 ));
    InMux I__3022 (
            .O(N__15088),
            .I(N__15082));
    InMux I__3021 (
            .O(N__15087),
            .I(N__15082));
    LocalMux I__3020 (
            .O(N__15082),
            .I(N__15079));
    Odrv12 I__3019 (
            .O(N__15079),
            .I(\Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ));
    InMux I__3018 (
            .O(N__15076),
            .I(N__15073));
    LocalMux I__3017 (
            .O(N__15073),
            .I(\Lab_UT.dictrl.g0_3_4 ));
    InMux I__3016 (
            .O(N__15070),
            .I(N__15067));
    LocalMux I__3015 (
            .O(N__15067),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0 ));
    InMux I__3014 (
            .O(N__15064),
            .I(N__15061));
    LocalMux I__3013 (
            .O(N__15061),
            .I(N__15058));
    Odrv4 I__3012 (
            .O(N__15058),
            .I(\Lab_UT.dictrl.G_14_0_a2_4_2 ));
    CascadeMux I__3011 (
            .O(N__15055),
            .I(N__15051));
    CascadeMux I__3010 (
            .O(N__15054),
            .I(N__15048));
    InMux I__3009 (
            .O(N__15051),
            .I(N__15037));
    InMux I__3008 (
            .O(N__15048),
            .I(N__15037));
    InMux I__3007 (
            .O(N__15047),
            .I(N__15037));
    InMux I__3006 (
            .O(N__15046),
            .I(N__15037));
    LocalMux I__3005 (
            .O(N__15037),
            .I(N__15034));
    Odrv4 I__3004 (
            .O(N__15034),
            .I(\Lab_UT.dictrl.G_14_0_0 ));
    CascadeMux I__3003 (
            .O(N__15031),
            .I(N__15028));
    InMux I__3002 (
            .O(N__15028),
            .I(N__15025));
    LocalMux I__3001 (
            .O(N__15025),
            .I(\Lab_UT.dictrl.g2_0_0 ));
    CascadeMux I__3000 (
            .O(N__15022),
            .I(N__15019));
    InMux I__2999 (
            .O(N__15019),
            .I(N__15016));
    LocalMux I__2998 (
            .O(N__15016),
            .I(shifter_1_rep1_RNI0FPF));
    CascadeMux I__2997 (
            .O(N__15013),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ));
    InMux I__2996 (
            .O(N__15010),
            .I(N__14998));
    InMux I__2995 (
            .O(N__15009),
            .I(N__14998));
    InMux I__2994 (
            .O(N__15008),
            .I(N__14998));
    InMux I__2993 (
            .O(N__15007),
            .I(N__14998));
    LocalMux I__2992 (
            .O(N__14998),
            .I(N__14995));
    Odrv4 I__2991 (
            .O(N__14995),
            .I(\Lab_UT.dictrl.G_14_0_1 ));
    InMux I__2990 (
            .O(N__14992),
            .I(N__14989));
    LocalMux I__2989 (
            .O(N__14989),
            .I(N_15));
    CascadeMux I__2988 (
            .O(N__14986),
            .I(\Lab_UT.dictrl.G_14_0_a2_1_cascade_ ));
    InMux I__2987 (
            .O(N__14983),
            .I(N__14977));
    InMux I__2986 (
            .O(N__14982),
            .I(N__14977));
    LocalMux I__2985 (
            .O(N__14977),
            .I(N_14_0));
    CascadeMux I__2984 (
            .O(N__14974),
            .I(N__14968));
    CascadeMux I__2983 (
            .O(N__14973),
            .I(N__14965));
    InMux I__2982 (
            .O(N__14972),
            .I(N__14956));
    InMux I__2981 (
            .O(N__14971),
            .I(N__14956));
    InMux I__2980 (
            .O(N__14968),
            .I(N__14956));
    InMux I__2979 (
            .O(N__14965),
            .I(N__14956));
    LocalMux I__2978 (
            .O(N__14956),
            .I(N__14953));
    Span4Mux_h I__2977 (
            .O(N__14953),
            .I(N__14950));
    Odrv4 I__2976 (
            .O(N__14950),
            .I(\Lab_UT.dictrl.N_20_0 ));
    CascadeMux I__2975 (
            .O(N__14947),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_ ));
    InMux I__2974 (
            .O(N__14944),
            .I(N__14940));
    InMux I__2973 (
            .O(N__14943),
            .I(N__14937));
    LocalMux I__2972 (
            .O(N__14940),
            .I(\Lab_UT.dictrl.N_22 ));
    LocalMux I__2971 (
            .O(N__14937),
            .I(\Lab_UT.dictrl.N_22 ));
    CascadeMux I__2970 (
            .O(N__14932),
            .I(N__14929));
    InMux I__2969 (
            .O(N__14929),
            .I(N__14926));
    LocalMux I__2968 (
            .O(N__14926),
            .I(\Lab_UT.dictrl.next_state_0_1 ));
    CascadeMux I__2967 (
            .O(N__14923),
            .I(\Lab_UT.dictrl.N_20_0_0_cascade_ ));
    InMux I__2966 (
            .O(N__14920),
            .I(N__14917));
    LocalMux I__2965 (
            .O(N__14917),
            .I(\Lab_UT.dictrl.N_22_0_0 ));
    InMux I__2964 (
            .O(N__14914),
            .I(N__14911));
    LocalMux I__2963 (
            .O(N__14911),
            .I(\Lab_UT.didp.g0_0Z0Z_2 ));
    CascadeMux I__2962 (
            .O(N__14908),
            .I(\Lab_UT.next_state_1_0_0_1_cascade_ ));
    InMux I__2961 (
            .O(N__14905),
            .I(N__14899));
    InMux I__2960 (
            .O(N__14904),
            .I(N__14899));
    LocalMux I__2959 (
            .O(N__14899),
            .I(N__14896));
    Odrv4 I__2958 (
            .O(N__14896),
            .I(\Lab_UT.dictrl.next_state6 ));
    InMux I__2957 (
            .O(N__14893),
            .I(N__14887));
    InMux I__2956 (
            .O(N__14892),
            .I(N__14887));
    LocalMux I__2955 (
            .O(N__14887),
            .I(\Lab_UT.dictrl.m19_1 ));
    CascadeMux I__2954 (
            .O(N__14884),
            .I(N__14881));
    InMux I__2953 (
            .O(N__14881),
            .I(N__14878));
    LocalMux I__2952 (
            .O(N__14878),
            .I(N__14875));
    Odrv12 I__2951 (
            .O(N__14875),
            .I(\Lab_UT.dictrl.m19_1_0 ));
    InMux I__2950 (
            .O(N__14872),
            .I(N__14868));
    CascadeMux I__2949 (
            .O(N__14871),
            .I(N__14864));
    LocalMux I__2948 (
            .O(N__14868),
            .I(N__14861));
    InMux I__2947 (
            .O(N__14867),
            .I(N__14858));
    InMux I__2946 (
            .O(N__14864),
            .I(N__14855));
    Odrv4 I__2945 (
            .O(N__14861),
            .I(\Lab_UT.dictrl.N_20 ));
    LocalMux I__2944 (
            .O(N__14858),
            .I(\Lab_UT.dictrl.N_20 ));
    LocalMux I__2943 (
            .O(N__14855),
            .I(\Lab_UT.dictrl.N_20 ));
    InMux I__2942 (
            .O(N__14848),
            .I(N__14845));
    LocalMux I__2941 (
            .O(N__14845),
            .I(N__14840));
    InMux I__2940 (
            .O(N__14844),
            .I(N__14837));
    InMux I__2939 (
            .O(N__14843),
            .I(N__14834));
    Odrv4 I__2938 (
            .O(N__14840),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    LocalMux I__2937 (
            .O(N__14837),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    LocalMux I__2936 (
            .O(N__14834),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    CascadeMux I__2935 (
            .O(N__14827),
            .I(\Lab_UT.dictrl.N_20_cascade_ ));
    CascadeMux I__2934 (
            .O(N__14824),
            .I(N__14821));
    InMux I__2933 (
            .O(N__14821),
            .I(N__14817));
    InMux I__2932 (
            .O(N__14820),
            .I(N__14814));
    LocalMux I__2931 (
            .O(N__14817),
            .I(\Lab_UT.dictrl.dicRun_1 ));
    LocalMux I__2930 (
            .O(N__14814),
            .I(\Lab_UT.dictrl.dicRun_1 ));
    InMux I__2929 (
            .O(N__14809),
            .I(N__14805));
    InMux I__2928 (
            .O(N__14808),
            .I(N__14802));
    LocalMux I__2927 (
            .O(N__14805),
            .I(\Lab_UT.LdASones ));
    LocalMux I__2926 (
            .O(N__14802),
            .I(\Lab_UT.LdASones ));
    InMux I__2925 (
            .O(N__14797),
            .I(N__14794));
    LocalMux I__2924 (
            .O(N__14794),
            .I(N__14791));
    Span4Mux_s3_h I__2923 (
            .O(N__14791),
            .I(N__14787));
    InMux I__2922 (
            .O(N__14790),
            .I(N__14784));
    Span4Mux_h I__2921 (
            .O(N__14787),
            .I(N__14781));
    LocalMux I__2920 (
            .O(N__14784),
            .I(N__14778));
    Odrv4 I__2919 (
            .O(N__14781),
            .I(\Lab_UT.LdAStens ));
    Odrv4 I__2918 (
            .O(N__14778),
            .I(\Lab_UT.LdAStens ));
    InMux I__2917 (
            .O(N__14773),
            .I(N__14764));
    InMux I__2916 (
            .O(N__14772),
            .I(N__14764));
    InMux I__2915 (
            .O(N__14771),
            .I(N__14764));
    LocalMux I__2914 (
            .O(N__14764),
            .I(N__14761));
    Span4Mux_v I__2913 (
            .O(N__14761),
            .I(N__14758));
    Odrv4 I__2912 (
            .O(N__14758),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    CascadeMux I__2911 (
            .O(N__14755),
            .I(N__14751));
    CascadeMux I__2910 (
            .O(N__14754),
            .I(N__14748));
    InMux I__2909 (
            .O(N__14751),
            .I(N__14743));
    InMux I__2908 (
            .O(N__14748),
            .I(N__14738));
    InMux I__2907 (
            .O(N__14747),
            .I(N__14738));
    InMux I__2906 (
            .O(N__14746),
            .I(N__14735));
    LocalMux I__2905 (
            .O(N__14743),
            .I(N__14732));
    LocalMux I__2904 (
            .O(N__14738),
            .I(N__14729));
    LocalMux I__2903 (
            .O(N__14735),
            .I(N__14726));
    Span4Mux_h I__2902 (
            .O(N__14732),
            .I(N__14721));
    Span4Mux_h I__2901 (
            .O(N__14729),
            .I(N__14721));
    Span4Mux_h I__2900 (
            .O(N__14726),
            .I(N__14718));
    Odrv4 I__2899 (
            .O(N__14721),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    Odrv4 I__2898 (
            .O(N__14718),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    InMux I__2897 (
            .O(N__14713),
            .I(N__14707));
    InMux I__2896 (
            .O(N__14712),
            .I(N__14707));
    LocalMux I__2895 (
            .O(N__14707),
            .I(\Lab_UT.dictrl.dicLdAMones_1 ));
    InMux I__2894 (
            .O(N__14704),
            .I(N__14701));
    LocalMux I__2893 (
            .O(N__14701),
            .I(N__14698));
    Span4Mux_h I__2892 (
            .O(N__14698),
            .I(N__14695));
    Odrv4 I__2891 (
            .O(N__14695),
            .I(\Lab_UT.LdAMones ));
    CascadeMux I__2890 (
            .O(N__14692),
            .I(\Lab_UT.LdAMones_cascade_ ));
    InMux I__2889 (
            .O(N__14689),
            .I(N__14686));
    LocalMux I__2888 (
            .O(N__14686),
            .I(N__14683));
    Span4Mux_h I__2887 (
            .O(N__14683),
            .I(N__14680));
    Span4Mux_v I__2886 (
            .O(N__14680),
            .I(N__14677));
    Odrv4 I__2885 (
            .O(N__14677),
            .I(\Lab_UT.dictrl.state_ret_2_fast ));
    InMux I__2884 (
            .O(N__14674),
            .I(N__14671));
    LocalMux I__2883 (
            .O(N__14671),
            .I(\uu2.bitmapZ0Z_72 ));
    InMux I__2882 (
            .O(N__14668),
            .I(N__14659));
    InMux I__2881 (
            .O(N__14667),
            .I(N__14659));
    InMux I__2880 (
            .O(N__14666),
            .I(N__14659));
    LocalMux I__2879 (
            .O(N__14659),
            .I(N__14654));
    InMux I__2878 (
            .O(N__14658),
            .I(N__14649));
    InMux I__2877 (
            .O(N__14657),
            .I(N__14649));
    Span4Mux_s1_v I__2876 (
            .O(N__14654),
            .I(N__14644));
    LocalMux I__2875 (
            .O(N__14649),
            .I(N__14641));
    InMux I__2874 (
            .O(N__14648),
            .I(N__14636));
    InMux I__2873 (
            .O(N__14647),
            .I(N__14636));
    Odrv4 I__2872 (
            .O(N__14644),
            .I(\Lab_UT.min2_2 ));
    Odrv4 I__2871 (
            .O(N__14641),
            .I(\Lab_UT.min2_2 ));
    LocalMux I__2870 (
            .O(N__14636),
            .I(\Lab_UT.min2_2 ));
    CascadeMux I__2869 (
            .O(N__14629),
            .I(N__14623));
    CascadeMux I__2868 (
            .O(N__14628),
            .I(N__14618));
    CascadeMux I__2867 (
            .O(N__14627),
            .I(N__14615));
    InMux I__2866 (
            .O(N__14626),
            .I(N__14610));
    InMux I__2865 (
            .O(N__14623),
            .I(N__14610));
    CascadeMux I__2864 (
            .O(N__14622),
            .I(N__14606));
    InMux I__2863 (
            .O(N__14621),
            .I(N__14599));
    InMux I__2862 (
            .O(N__14618),
            .I(N__14599));
    InMux I__2861 (
            .O(N__14615),
            .I(N__14599));
    LocalMux I__2860 (
            .O(N__14610),
            .I(N__14596));
    InMux I__2859 (
            .O(N__14609),
            .I(N__14591));
    InMux I__2858 (
            .O(N__14606),
            .I(N__14591));
    LocalMux I__2857 (
            .O(N__14599),
            .I(\Lab_UT.min2_3 ));
    Odrv12 I__2856 (
            .O(N__14596),
            .I(\Lab_UT.min2_3 ));
    LocalMux I__2855 (
            .O(N__14591),
            .I(\Lab_UT.min2_3 ));
    InMux I__2854 (
            .O(N__14584),
            .I(N__14578));
    InMux I__2853 (
            .O(N__14583),
            .I(N__14578));
    LocalMux I__2852 (
            .O(N__14578),
            .I(N__14572));
    InMux I__2851 (
            .O(N__14577),
            .I(N__14565));
    InMux I__2850 (
            .O(N__14576),
            .I(N__14565));
    InMux I__2849 (
            .O(N__14575),
            .I(N__14565));
    Span4Mux_s3_v I__2848 (
            .O(N__14572),
            .I(N__14560));
    LocalMux I__2847 (
            .O(N__14565),
            .I(N__14557));
    InMux I__2846 (
            .O(N__14564),
            .I(N__14552));
    InMux I__2845 (
            .O(N__14563),
            .I(N__14552));
    Odrv4 I__2844 (
            .O(N__14560),
            .I(\Lab_UT.min2_0 ));
    Odrv12 I__2843 (
            .O(N__14557),
            .I(\Lab_UT.min2_0 ));
    LocalMux I__2842 (
            .O(N__14552),
            .I(\Lab_UT.min2_0 ));
    CascadeMux I__2841 (
            .O(N__14545),
            .I(N__14542));
    InMux I__2840 (
            .O(N__14542),
            .I(N__14539));
    LocalMux I__2839 (
            .O(N__14539),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__2838 (
            .O(N__14536),
            .I(N__14533));
    LocalMux I__2837 (
            .O(N__14533),
            .I(N__14528));
    InMux I__2836 (
            .O(N__14532),
            .I(N__14525));
    InMux I__2835 (
            .O(N__14531),
            .I(N__14522));
    Span4Mux_h I__2834 (
            .O(N__14528),
            .I(N__14517));
    LocalMux I__2833 (
            .O(N__14525),
            .I(N__14517));
    LocalMux I__2832 (
            .O(N__14522),
            .I(N__14514));
    Span4Mux_h I__2831 (
            .O(N__14517),
            .I(N__14511));
    Odrv4 I__2830 (
            .O(N__14514),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__2829 (
            .O(N__14511),
            .I(\Lab_UT.di_AMones_1 ));
    CascadeMux I__2828 (
            .O(N__14506),
            .I(N__14503));
    InMux I__2827 (
            .O(N__14503),
            .I(N__14492));
    InMux I__2826 (
            .O(N__14502),
            .I(N__14492));
    InMux I__2825 (
            .O(N__14501),
            .I(N__14492));
    CascadeMux I__2824 (
            .O(N__14500),
            .I(N__14489));
    CascadeMux I__2823 (
            .O(N__14499),
            .I(N__14485));
    LocalMux I__2822 (
            .O(N__14492),
            .I(N__14481));
    InMux I__2821 (
            .O(N__14489),
            .I(N__14476));
    InMux I__2820 (
            .O(N__14488),
            .I(N__14476));
    InMux I__2819 (
            .O(N__14485),
            .I(N__14471));
    InMux I__2818 (
            .O(N__14484),
            .I(N__14471));
    Span4Mux_s1_v I__2817 (
            .O(N__14481),
            .I(N__14468));
    LocalMux I__2816 (
            .O(N__14476),
            .I(N__14465));
    LocalMux I__2815 (
            .O(N__14471),
            .I(N__14462));
    Odrv4 I__2814 (
            .O(N__14468),
            .I(\Lab_UT.min2_1 ));
    Odrv12 I__2813 (
            .O(N__14465),
            .I(\Lab_UT.min2_1 ));
    Odrv4 I__2812 (
            .O(N__14462),
            .I(\Lab_UT.min2_1 ));
    CascadeMux I__2811 (
            .O(N__14455),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__2810 (
            .O(N__14452),
            .I(N__14445));
    InMux I__2809 (
            .O(N__14451),
            .I(N__14445));
    InMux I__2808 (
            .O(N__14450),
            .I(N__14442));
    LocalMux I__2807 (
            .O(N__14445),
            .I(N__14439));
    LocalMux I__2806 (
            .O(N__14442),
            .I(N__14434));
    Span4Mux_h I__2805 (
            .O(N__14439),
            .I(N__14429));
    InMux I__2804 (
            .O(N__14438),
            .I(N__14426));
    InMux I__2803 (
            .O(N__14437),
            .I(N__14423));
    Span4Mux_v I__2802 (
            .O(N__14434),
            .I(N__14420));
    InMux I__2801 (
            .O(N__14433),
            .I(N__14415));
    InMux I__2800 (
            .O(N__14432),
            .I(N__14415));
    Span4Mux_s2_v I__2799 (
            .O(N__14429),
            .I(N__14412));
    LocalMux I__2798 (
            .O(N__14426),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__2797 (
            .O(N__14423),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__2796 (
            .O(N__14420),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__2795 (
            .O(N__14415),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__2794 (
            .O(N__14412),
            .I(\Lab_UT.di_Mtens_0 ));
    InMux I__2793 (
            .O(N__14401),
            .I(N__14397));
    InMux I__2792 (
            .O(N__14400),
            .I(N__14393));
    LocalMux I__2791 (
            .O(N__14397),
            .I(N__14390));
    InMux I__2790 (
            .O(N__14396),
            .I(N__14387));
    LocalMux I__2789 (
            .O(N__14393),
            .I(N__14384));
    Span4Mux_v I__2788 (
            .O(N__14390),
            .I(N__14379));
    LocalMux I__2787 (
            .O(N__14387),
            .I(N__14379));
    Odrv4 I__2786 (
            .O(N__14384),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__2785 (
            .O(N__14379),
            .I(\Lab_UT.di_ASones_2 ));
    InMux I__2784 (
            .O(N__14374),
            .I(N__14371));
    LocalMux I__2783 (
            .O(N__14371),
            .I(N__14368));
    Span4Mux_h I__2782 (
            .O(N__14368),
            .I(N__14365));
    Odrv4 I__2781 (
            .O(N__14365),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ));
    InMux I__2780 (
            .O(N__14362),
            .I(N__14359));
    LocalMux I__2779 (
            .O(N__14359),
            .I(N__14354));
    InMux I__2778 (
            .O(N__14358),
            .I(N__14351));
    InMux I__2777 (
            .O(N__14357),
            .I(N__14348));
    Span4Mux_h I__2776 (
            .O(N__14354),
            .I(N__14344));
    LocalMux I__2775 (
            .O(N__14351),
            .I(N__14339));
    LocalMux I__2774 (
            .O(N__14348),
            .I(N__14339));
    InMux I__2773 (
            .O(N__14347),
            .I(N__14336));
    Span4Mux_h I__2772 (
            .O(N__14344),
            .I(N__14333));
    Odrv12 I__2771 (
            .O(N__14339),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__2770 (
            .O(N__14336),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__2769 (
            .O(N__14333),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__2768 (
            .O(N__14326),
            .I(N__14323));
    LocalMux I__2767 (
            .O(N__14323),
            .I(N__14319));
    InMux I__2766 (
            .O(N__14322),
            .I(N__14316));
    Span4Mux_h I__2765 (
            .O(N__14319),
            .I(N__14311));
    LocalMux I__2764 (
            .O(N__14316),
            .I(N__14311));
    Span4Mux_h I__2763 (
            .O(N__14311),
            .I(N__14308));
    Odrv4 I__2762 (
            .O(N__14308),
            .I(\uu2.un1_l_count_1_0 ));
    CascadeMux I__2761 (
            .O(N__14305),
            .I(N__14302));
    InMux I__2760 (
            .O(N__14302),
            .I(N__14293));
    InMux I__2759 (
            .O(N__14301),
            .I(N__14290));
    InMux I__2758 (
            .O(N__14300),
            .I(N__14285));
    InMux I__2757 (
            .O(N__14299),
            .I(N__14285));
    InMux I__2756 (
            .O(N__14298),
            .I(N__14278));
    InMux I__2755 (
            .O(N__14297),
            .I(N__14278));
    InMux I__2754 (
            .O(N__14296),
            .I(N__14278));
    LocalMux I__2753 (
            .O(N__14293),
            .I(N__14275));
    LocalMux I__2752 (
            .O(N__14290),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2751 (
            .O(N__14285),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2750 (
            .O(N__14278),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv12 I__2749 (
            .O(N__14275),
            .I(\Lab_UT.di_Stens_0 ));
    InMux I__2748 (
            .O(N__14266),
            .I(N__14261));
    InMux I__2747 (
            .O(N__14265),
            .I(N__14254));
    InMux I__2746 (
            .O(N__14264),
            .I(N__14250));
    LocalMux I__2745 (
            .O(N__14261),
            .I(N__14247));
    InMux I__2744 (
            .O(N__14260),
            .I(N__14244));
    InMux I__2743 (
            .O(N__14259),
            .I(N__14241));
    InMux I__2742 (
            .O(N__14258),
            .I(N__14238));
    InMux I__2741 (
            .O(N__14257),
            .I(N__14235));
    LocalMux I__2740 (
            .O(N__14254),
            .I(N__14232));
    InMux I__2739 (
            .O(N__14253),
            .I(N__14229));
    LocalMux I__2738 (
            .O(N__14250),
            .I(N__14224));
    Span4Mux_h I__2737 (
            .O(N__14247),
            .I(N__14224));
    LocalMux I__2736 (
            .O(N__14244),
            .I(N__14216));
    LocalMux I__2735 (
            .O(N__14241),
            .I(N__14211));
    LocalMux I__2734 (
            .O(N__14238),
            .I(N__14211));
    LocalMux I__2733 (
            .O(N__14235),
            .I(N__14206));
    Span4Mux_v I__2732 (
            .O(N__14232),
            .I(N__14206));
    LocalMux I__2731 (
            .O(N__14229),
            .I(N__14201));
    Span4Mux_v I__2730 (
            .O(N__14224),
            .I(N__14201));
    InMux I__2729 (
            .O(N__14223),
            .I(N__14196));
    InMux I__2728 (
            .O(N__14222),
            .I(N__14196));
    InMux I__2727 (
            .O(N__14221),
            .I(N__14189));
    InMux I__2726 (
            .O(N__14220),
            .I(N__14189));
    InMux I__2725 (
            .O(N__14219),
            .I(N__14189));
    Span4Mux_v I__2724 (
            .O(N__14216),
            .I(N__14186));
    Span4Mux_v I__2723 (
            .O(N__14211),
            .I(N__14183));
    Span4Mux_v I__2722 (
            .O(N__14206),
            .I(N__14178));
    Span4Mux_v I__2721 (
            .O(N__14201),
            .I(N__14178));
    LocalMux I__2720 (
            .O(N__14196),
            .I(N__14173));
    LocalMux I__2719 (
            .O(N__14189),
            .I(N__14173));
    Odrv4 I__2718 (
            .O(N__14186),
            .I(bu_rx_data_0));
    Odrv4 I__2717 (
            .O(N__14183),
            .I(bu_rx_data_0));
    Odrv4 I__2716 (
            .O(N__14178),
            .I(bu_rx_data_0));
    Odrv12 I__2715 (
            .O(N__14173),
            .I(bu_rx_data_0));
    InMux I__2714 (
            .O(N__14164),
            .I(N__14161));
    LocalMux I__2713 (
            .O(N__14161),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ));
    InMux I__2712 (
            .O(N__14158),
            .I(N__14155));
    LocalMux I__2711 (
            .O(N__14155),
            .I(N__14150));
    InMux I__2710 (
            .O(N__14154),
            .I(N__14147));
    InMux I__2709 (
            .O(N__14153),
            .I(N__14144));
    Span4Mux_v I__2708 (
            .O(N__14150),
            .I(N__14139));
    LocalMux I__2707 (
            .O(N__14147),
            .I(N__14139));
    LocalMux I__2706 (
            .O(N__14144),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__2705 (
            .O(N__14139),
            .I(\Lab_UT.di_AMones_2 ));
    CascadeMux I__2704 (
            .O(N__14134),
            .I(N__14127));
    CascadeMux I__2703 (
            .O(N__14133),
            .I(N__14124));
    CascadeMux I__2702 (
            .O(N__14132),
            .I(N__14121));
    CascadeMux I__2701 (
            .O(N__14131),
            .I(N__14118));
    InMux I__2700 (
            .O(N__14130),
            .I(N__14113));
    InMux I__2699 (
            .O(N__14127),
            .I(N__14100));
    InMux I__2698 (
            .O(N__14124),
            .I(N__14100));
    InMux I__2697 (
            .O(N__14121),
            .I(N__14100));
    InMux I__2696 (
            .O(N__14118),
            .I(N__14100));
    InMux I__2695 (
            .O(N__14117),
            .I(N__14100));
    InMux I__2694 (
            .O(N__14116),
            .I(N__14100));
    LocalMux I__2693 (
            .O(N__14113),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__2692 (
            .O(N__14100),
            .I(\Lab_UT.sec1_1 ));
    InMux I__2691 (
            .O(N__14095),
            .I(N__14086));
    InMux I__2690 (
            .O(N__14094),
            .I(N__14073));
    InMux I__2689 (
            .O(N__14093),
            .I(N__14073));
    InMux I__2688 (
            .O(N__14092),
            .I(N__14073));
    InMux I__2687 (
            .O(N__14091),
            .I(N__14073));
    InMux I__2686 (
            .O(N__14090),
            .I(N__14073));
    InMux I__2685 (
            .O(N__14089),
            .I(N__14073));
    LocalMux I__2684 (
            .O(N__14086),
            .I(\Lab_UT.sec1_2 ));
    LocalMux I__2683 (
            .O(N__14073),
            .I(\Lab_UT.sec1_2 ));
    CascadeMux I__2682 (
            .O(N__14068),
            .I(N__14059));
    CascadeMux I__2681 (
            .O(N__14067),
            .I(N__14056));
    CascadeMux I__2680 (
            .O(N__14066),
            .I(N__14053));
    InMux I__2679 (
            .O(N__14065),
            .I(N__14040));
    InMux I__2678 (
            .O(N__14064),
            .I(N__14040));
    InMux I__2677 (
            .O(N__14063),
            .I(N__14040));
    InMux I__2676 (
            .O(N__14062),
            .I(N__14040));
    InMux I__2675 (
            .O(N__14059),
            .I(N__14040));
    InMux I__2674 (
            .O(N__14056),
            .I(N__14040));
    InMux I__2673 (
            .O(N__14053),
            .I(N__14037));
    LocalMux I__2672 (
            .O(N__14040),
            .I(N__14034));
    LocalMux I__2671 (
            .O(N__14037),
            .I(\Lab_UT.sec1_3 ));
    Odrv4 I__2670 (
            .O(N__14034),
            .I(\Lab_UT.sec1_3 ));
    InMux I__2669 (
            .O(N__14029),
            .I(N__14020));
    InMux I__2668 (
            .O(N__14028),
            .I(N__14007));
    InMux I__2667 (
            .O(N__14027),
            .I(N__14007));
    InMux I__2666 (
            .O(N__14026),
            .I(N__14007));
    InMux I__2665 (
            .O(N__14025),
            .I(N__14007));
    InMux I__2664 (
            .O(N__14024),
            .I(N__14007));
    InMux I__2663 (
            .O(N__14023),
            .I(N__14007));
    LocalMux I__2662 (
            .O(N__14020),
            .I(\Lab_UT.sec1_0 ));
    LocalMux I__2661 (
            .O(N__14007),
            .I(\Lab_UT.sec1_0 ));
    InMux I__2660 (
            .O(N__14002),
            .I(N__13999));
    LocalMux I__2659 (
            .O(N__13999),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__2658 (
            .O(N__13996),
            .I(N__13993));
    LocalMux I__2657 (
            .O(N__13993),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__2656 (
            .O(N__13990),
            .I(N__13987));
    LocalMux I__2655 (
            .O(N__13987),
            .I(\uu2.bitmap_pmux_17_ns_1 ));
    CascadeMux I__2654 (
            .O(N__13984),
            .I(N__13979));
    InMux I__2653 (
            .O(N__13983),
            .I(N__13972));
    InMux I__2652 (
            .O(N__13982),
            .I(N__13972));
    InMux I__2651 (
            .O(N__13979),
            .I(N__13972));
    LocalMux I__2650 (
            .O(N__13972),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__2649 (
            .O(N__13969),
            .I(N__13966));
    LocalMux I__2648 (
            .O(N__13966),
            .I(N__13963));
    Odrv4 I__2647 (
            .O(N__13963),
            .I(\uu2.bitmap_pmux_16_ns_1 ));
    CascadeMux I__2646 (
            .O(N__13960),
            .I(N__13954));
    InMux I__2645 (
            .O(N__13959),
            .I(N__13948));
    InMux I__2644 (
            .O(N__13958),
            .I(N__13948));
    InMux I__2643 (
            .O(N__13957),
            .I(N__13936));
    InMux I__2642 (
            .O(N__13954),
            .I(N__13936));
    InMux I__2641 (
            .O(N__13953),
            .I(N__13936));
    LocalMux I__2640 (
            .O(N__13948),
            .I(N__13933));
    InMux I__2639 (
            .O(N__13947),
            .I(N__13925));
    InMux I__2638 (
            .O(N__13946),
            .I(N__13925));
    InMux I__2637 (
            .O(N__13945),
            .I(N__13925));
    InMux I__2636 (
            .O(N__13944),
            .I(N__13920));
    InMux I__2635 (
            .O(N__13943),
            .I(N__13920));
    LocalMux I__2634 (
            .O(N__13936),
            .I(N__13917));
    Span4Mux_v I__2633 (
            .O(N__13933),
            .I(N__13914));
    InMux I__2632 (
            .O(N__13932),
            .I(N__13911));
    LocalMux I__2631 (
            .O(N__13925),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    LocalMux I__2630 (
            .O(N__13920),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    Odrv4 I__2629 (
            .O(N__13917),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    Odrv4 I__2628 (
            .O(N__13914),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    LocalMux I__2627 (
            .O(N__13911),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    InMux I__2626 (
            .O(N__13900),
            .I(N__13897));
    LocalMux I__2625 (
            .O(N__13897),
            .I(N__13893));
    InMux I__2624 (
            .O(N__13896),
            .I(N__13890));
    Span4Mux_v I__2623 (
            .O(N__13893),
            .I(N__13885));
    LocalMux I__2622 (
            .O(N__13890),
            .I(N__13885));
    Span4Mux_h I__2621 (
            .O(N__13885),
            .I(N__13882));
    Odrv4 I__2620 (
            .O(N__13882),
            .I(\uu2.N_44 ));
    CascadeMux I__2619 (
            .O(N__13879),
            .I(N__13875));
    InMux I__2618 (
            .O(N__13878),
            .I(N__13872));
    InMux I__2617 (
            .O(N__13875),
            .I(N__13868));
    LocalMux I__2616 (
            .O(N__13872),
            .I(N__13865));
    InMux I__2615 (
            .O(N__13871),
            .I(N__13862));
    LocalMux I__2614 (
            .O(N__13868),
            .I(N__13859));
    Span4Mux_h I__2613 (
            .O(N__13865),
            .I(N__13856));
    LocalMux I__2612 (
            .O(N__13862),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__2611 (
            .O(N__13859),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__2610 (
            .O(N__13856),
            .I(\Lab_UT.di_AMtens_0 ));
    InMux I__2609 (
            .O(N__13849),
            .I(N__13846));
    LocalMux I__2608 (
            .O(N__13846),
            .I(N__13843));
    Span4Mux_v I__2607 (
            .O(N__13843),
            .I(N__13840));
    Odrv4 I__2606 (
            .O(N__13840),
            .I(\Lab_UT.didp.reset_12_1_3 ));
    InMux I__2605 (
            .O(N__13837),
            .I(N__13834));
    LocalMux I__2604 (
            .O(N__13834),
            .I(N__13831));
    Span4Mux_v I__2603 (
            .O(N__13831),
            .I(N__13828));
    Span4Mux_h I__2602 (
            .O(N__13828),
            .I(N__13823));
    InMux I__2601 (
            .O(N__13827),
            .I(N__13818));
    InMux I__2600 (
            .O(N__13826),
            .I(N__13818));
    Odrv4 I__2599 (
            .O(N__13823),
            .I(\Lab_UT.di_AMtens_3 ));
    LocalMux I__2598 (
            .O(N__13818),
            .I(\Lab_UT.di_AMtens_3 ));
    InMux I__2597 (
            .O(N__13813),
            .I(N__13810));
    LocalMux I__2596 (
            .O(N__13810),
            .I(N__13806));
    InMux I__2595 (
            .O(N__13809),
            .I(N__13803));
    Span4Mux_s3_v I__2594 (
            .O(N__13806),
            .I(N__13800));
    LocalMux I__2593 (
            .O(N__13803),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__2592 (
            .O(N__13800),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__2591 (
            .O(N__13795),
            .I(N__13792));
    LocalMux I__2590 (
            .O(N__13792),
            .I(N__13789));
    Span4Mux_h I__2589 (
            .O(N__13789),
            .I(N__13786));
    Span4Mux_v I__2588 (
            .O(N__13786),
            .I(N__13781));
    InMux I__2587 (
            .O(N__13785),
            .I(N__13778));
    InMux I__2586 (
            .O(N__13784),
            .I(N__13775));
    Span4Mux_h I__2585 (
            .O(N__13781),
            .I(N__13772));
    LocalMux I__2584 (
            .O(N__13778),
            .I(\buart.Z_rx.idle ));
    LocalMux I__2583 (
            .O(N__13775),
            .I(\buart.Z_rx.idle ));
    Odrv4 I__2582 (
            .O(N__13772),
            .I(\buart.Z_rx.idle ));
    InMux I__2581 (
            .O(N__13765),
            .I(N__13761));
    CascadeMux I__2580 (
            .O(N__13764),
            .I(N__13754));
    LocalMux I__2579 (
            .O(N__13761),
            .I(N__13745));
    InMux I__2578 (
            .O(N__13760),
            .I(N__13742));
    InMux I__2577 (
            .O(N__13759),
            .I(N__13739));
    InMux I__2576 (
            .O(N__13758),
            .I(N__13736));
    InMux I__2575 (
            .O(N__13757),
            .I(N__13733));
    InMux I__2574 (
            .O(N__13754),
            .I(N__13730));
    InMux I__2573 (
            .O(N__13753),
            .I(N__13721));
    InMux I__2572 (
            .O(N__13752),
            .I(N__13721));
    InMux I__2571 (
            .O(N__13751),
            .I(N__13721));
    InMux I__2570 (
            .O(N__13750),
            .I(N__13721));
    InMux I__2569 (
            .O(N__13749),
            .I(N__13716));
    InMux I__2568 (
            .O(N__13748),
            .I(N__13716));
    Span4Mux_v I__2567 (
            .O(N__13745),
            .I(N__13713));
    LocalMux I__2566 (
            .O(N__13742),
            .I(N__13706));
    LocalMux I__2565 (
            .O(N__13739),
            .I(N__13706));
    LocalMux I__2564 (
            .O(N__13736),
            .I(N__13706));
    LocalMux I__2563 (
            .O(N__13733),
            .I(N__13703));
    LocalMux I__2562 (
            .O(N__13730),
            .I(N__13698));
    LocalMux I__2561 (
            .O(N__13721),
            .I(N__13698));
    LocalMux I__2560 (
            .O(N__13716),
            .I(N__13691));
    Span4Mux_s1_h I__2559 (
            .O(N__13713),
            .I(N__13691));
    Span4Mux_v I__2558 (
            .O(N__13706),
            .I(N__13691));
    Span4Mux_h I__2557 (
            .O(N__13703),
            .I(N__13686));
    Span4Mux_h I__2556 (
            .O(N__13698),
            .I(N__13686));
    Sp12to4 I__2555 (
            .O(N__13691),
            .I(N__13683));
    Sp12to4 I__2554 (
            .O(N__13686),
            .I(N__13680));
    Span12Mux_s7_h I__2553 (
            .O(N__13683),
            .I(N__13677));
    Span12Mux_v I__2552 (
            .O(N__13680),
            .I(N__13674));
    Odrv12 I__2551 (
            .O(N__13677),
            .I(\buart.Z_rx.startbit ));
    Odrv12 I__2550 (
            .O(N__13674),
            .I(\buart.Z_rx.startbit ));
    InMux I__2549 (
            .O(N__13669),
            .I(N__13666));
    LocalMux I__2548 (
            .O(N__13666),
            .I(N__13663));
    Span4Mux_v I__2547 (
            .O(N__13663),
            .I(N__13658));
    InMux I__2546 (
            .O(N__13662),
            .I(N__13655));
    InMux I__2545 (
            .O(N__13661),
            .I(N__13652));
    Span4Mux_v I__2544 (
            .O(N__13658),
            .I(N__13649));
    LocalMux I__2543 (
            .O(N__13655),
            .I(N__13646));
    LocalMux I__2542 (
            .O(N__13652),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__2541 (
            .O(N__13649),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__2540 (
            .O(N__13646),
            .I(\Lab_UT.di_AStens_1 ));
    InMux I__2539 (
            .O(N__13639),
            .I(N__13635));
    InMux I__2538 (
            .O(N__13638),
            .I(N__13632));
    LocalMux I__2537 (
            .O(N__13635),
            .I(N__13628));
    LocalMux I__2536 (
            .O(N__13632),
            .I(N__13625));
    InMux I__2535 (
            .O(N__13631),
            .I(N__13622));
    Span4Mux_v I__2534 (
            .O(N__13628),
            .I(N__13619));
    Span4Mux_h I__2533 (
            .O(N__13625),
            .I(N__13614));
    LocalMux I__2532 (
            .O(N__13622),
            .I(N__13614));
    Odrv4 I__2531 (
            .O(N__13619),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__2530 (
            .O(N__13614),
            .I(\Lab_UT.di_ASones_1 ));
    CascadeMux I__2529 (
            .O(N__13609),
            .I(N__13603));
    InMux I__2528 (
            .O(N__13608),
            .I(N__13596));
    InMux I__2527 (
            .O(N__13607),
            .I(N__13596));
    InMux I__2526 (
            .O(N__13606),
            .I(N__13590));
    InMux I__2525 (
            .O(N__13603),
            .I(N__13590));
    InMux I__2524 (
            .O(N__13602),
            .I(N__13585));
    InMux I__2523 (
            .O(N__13601),
            .I(N__13585));
    LocalMux I__2522 (
            .O(N__13596),
            .I(N__13582));
    InMux I__2521 (
            .O(N__13595),
            .I(N__13579));
    LocalMux I__2520 (
            .O(N__13590),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__2519 (
            .O(N__13585),
            .I(\Lab_UT.di_Stens_1 ));
    Odrv4 I__2518 (
            .O(N__13582),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__2517 (
            .O(N__13579),
            .I(\Lab_UT.di_Stens_1 ));
    InMux I__2516 (
            .O(N__13570),
            .I(N__13567));
    LocalMux I__2515 (
            .O(N__13567),
            .I(\Lab_UT.didp.countrce2.N_93 ));
    InMux I__2514 (
            .O(N__13564),
            .I(N__13560));
    InMux I__2513 (
            .O(N__13563),
            .I(N__13555));
    LocalMux I__2512 (
            .O(N__13560),
            .I(N__13552));
    InMux I__2511 (
            .O(N__13559),
            .I(N__13547));
    InMux I__2510 (
            .O(N__13558),
            .I(N__13547));
    LocalMux I__2509 (
            .O(N__13555),
            .I(N__13543));
    Span4Mux_v I__2508 (
            .O(N__13552),
            .I(N__13538));
    LocalMux I__2507 (
            .O(N__13547),
            .I(N__13538));
    InMux I__2506 (
            .O(N__13546),
            .I(N__13535));
    Span12Mux_s3_v I__2505 (
            .O(N__13543),
            .I(N__13532));
    Span4Mux_h I__2504 (
            .O(N__13538),
            .I(N__13529));
    LocalMux I__2503 (
            .O(N__13535),
            .I(o_One_Sec_Pulse));
    Odrv12 I__2502 (
            .O(N__13532),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2501 (
            .O(N__13529),
            .I(o_One_Sec_Pulse));
    InMux I__2500 (
            .O(N__13522),
            .I(N__13519));
    LocalMux I__2499 (
            .O(N__13519),
            .I(\uu2.bitmapZ0Z_111 ));
    InMux I__2498 (
            .O(N__13516),
            .I(N__13513));
    LocalMux I__2497 (
            .O(N__13513),
            .I(N__13509));
    InMux I__2496 (
            .O(N__13512),
            .I(N__13506));
    Span4Mux_s1_v I__2495 (
            .O(N__13509),
            .I(N__13503));
    LocalMux I__2494 (
            .O(N__13506),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__2493 (
            .O(N__13503),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__2492 (
            .O(N__13498),
            .I(N__13495));
    LocalMux I__2491 (
            .O(N__13495),
            .I(N__13492));
    Span4Mux_s1_v I__2490 (
            .O(N__13492),
            .I(N__13489));
    Odrv4 I__2489 (
            .O(N__13489),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    CascadeMux I__2488 (
            .O(N__13486),
            .I(N__13483));
    InMux I__2487 (
            .O(N__13483),
            .I(N__13480));
    LocalMux I__2486 (
            .O(N__13480),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__2485 (
            .O(N__13477),
            .I(N__13474));
    LocalMux I__2484 (
            .O(N__13474),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__2483 (
            .O(N__13471),
            .I(N__13465));
    InMux I__2482 (
            .O(N__13470),
            .I(N__13455));
    InMux I__2481 (
            .O(N__13469),
            .I(N__13455));
    InMux I__2480 (
            .O(N__13468),
            .I(N__13455));
    LocalMux I__2479 (
            .O(N__13465),
            .I(N__13452));
    CascadeMux I__2478 (
            .O(N__13464),
            .I(N__13449));
    InMux I__2477 (
            .O(N__13463),
            .I(N__13446));
    InMux I__2476 (
            .O(N__13462),
            .I(N__13443));
    LocalMux I__2475 (
            .O(N__13455),
            .I(N__13438));
    Span4Mux_h I__2474 (
            .O(N__13452),
            .I(N__13438));
    InMux I__2473 (
            .O(N__13449),
            .I(N__13435));
    LocalMux I__2472 (
            .O(N__13446),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__2471 (
            .O(N__13443),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv4 I__2470 (
            .O(N__13438),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__2469 (
            .O(N__13435),
            .I(\Lab_UT.di_Sones_3 ));
    InMux I__2468 (
            .O(N__13426),
            .I(N__13421));
    InMux I__2467 (
            .O(N__13425),
            .I(N__13418));
    InMux I__2466 (
            .O(N__13424),
            .I(N__13415));
    LocalMux I__2465 (
            .O(N__13421),
            .I(N__13412));
    LocalMux I__2464 (
            .O(N__13418),
            .I(N__13409));
    LocalMux I__2463 (
            .O(N__13415),
            .I(N__13406));
    Span4Mux_v I__2462 (
            .O(N__13412),
            .I(N__13403));
    Span4Mux_h I__2461 (
            .O(N__13409),
            .I(N__13400));
    Odrv12 I__2460 (
            .O(N__13406),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__2459 (
            .O(N__13403),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__2458 (
            .O(N__13400),
            .I(\Lab_UT.di_ASones_3 ));
    InMux I__2457 (
            .O(N__13393),
            .I(N__13388));
    InMux I__2456 (
            .O(N__13392),
            .I(N__13383));
    InMux I__2455 (
            .O(N__13391),
            .I(N__13383));
    LocalMux I__2454 (
            .O(N__13388),
            .I(N__13380));
    LocalMux I__2453 (
            .O(N__13383),
            .I(N__13375));
    Span12Mux_s6_h I__2452 (
            .O(N__13380),
            .I(N__13375));
    Odrv12 I__2451 (
            .O(N__13375),
            .I(\Lab_UT.di_ASones_0 ));
    InMux I__2450 (
            .O(N__13372),
            .I(N__13368));
    InMux I__2449 (
            .O(N__13371),
            .I(N__13365));
    LocalMux I__2448 (
            .O(N__13368),
            .I(N__13362));
    LocalMux I__2447 (
            .O(N__13365),
            .I(N__13358));
    Span4Mux_v I__2446 (
            .O(N__13362),
            .I(N__13355));
    InMux I__2445 (
            .O(N__13361),
            .I(N__13352));
    Span4Mux_h I__2444 (
            .O(N__13358),
            .I(N__13349));
    Odrv4 I__2443 (
            .O(N__13355),
            .I(\Lab_UT.di_AMones_3 ));
    LocalMux I__2442 (
            .O(N__13352),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__2441 (
            .O(N__13349),
            .I(\Lab_UT.di_AMones_3 ));
    InMux I__2440 (
            .O(N__13342),
            .I(N__13333));
    InMux I__2439 (
            .O(N__13341),
            .I(N__13333));
    InMux I__2438 (
            .O(N__13340),
            .I(N__13330));
    InMux I__2437 (
            .O(N__13339),
            .I(N__13327));
    InMux I__2436 (
            .O(N__13338),
            .I(N__13322));
    LocalMux I__2435 (
            .O(N__13333),
            .I(N__13319));
    LocalMux I__2434 (
            .O(N__13330),
            .I(N__13316));
    LocalMux I__2433 (
            .O(N__13327),
            .I(N__13313));
    CascadeMux I__2432 (
            .O(N__13326),
            .I(N__13307));
    InMux I__2431 (
            .O(N__13325),
            .I(N__13304));
    LocalMux I__2430 (
            .O(N__13322),
            .I(N__13301));
    Span4Mux_h I__2429 (
            .O(N__13319),
            .I(N__13298));
    Span4Mux_h I__2428 (
            .O(N__13316),
            .I(N__13295));
    Span4Mux_h I__2427 (
            .O(N__13313),
            .I(N__13292));
    InMux I__2426 (
            .O(N__13312),
            .I(N__13283));
    InMux I__2425 (
            .O(N__13311),
            .I(N__13283));
    InMux I__2424 (
            .O(N__13310),
            .I(N__13283));
    InMux I__2423 (
            .O(N__13307),
            .I(N__13283));
    LocalMux I__2422 (
            .O(N__13304),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2421 (
            .O(N__13301),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2420 (
            .O(N__13298),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2419 (
            .O(N__13295),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2418 (
            .O(N__13292),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2417 (
            .O(N__13283),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CascadeMux I__2416 (
            .O(N__13270),
            .I(N__13267));
    InMux I__2415 (
            .O(N__13267),
            .I(N__13264));
    LocalMux I__2414 (
            .O(N__13264),
            .I(\uu2.N_45 ));
    CEMux I__2413 (
            .O(N__13261),
            .I(N__13257));
    CEMux I__2412 (
            .O(N__13260),
            .I(N__13254));
    LocalMux I__2411 (
            .O(N__13257),
            .I(N__13250));
    LocalMux I__2410 (
            .O(N__13254),
            .I(N__13247));
    CEMux I__2409 (
            .O(N__13253),
            .I(N__13244));
    Span4Mux_s3_v I__2408 (
            .O(N__13250),
            .I(N__13241));
    Span4Mux_s0_v I__2407 (
            .O(N__13247),
            .I(N__13238));
    LocalMux I__2406 (
            .O(N__13244),
            .I(N__13233));
    Span4Mux_h I__2405 (
            .O(N__13241),
            .I(N__13233));
    Odrv4 I__2404 (
            .O(N__13238),
            .I(\uu2.N_33_1 ));
    Odrv4 I__2403 (
            .O(N__13233),
            .I(\uu2.N_33_1 ));
    InMux I__2402 (
            .O(N__13228),
            .I(N__13225));
    LocalMux I__2401 (
            .O(N__13225),
            .I(N__13221));
    CascadeMux I__2400 (
            .O(N__13224),
            .I(N__13216));
    Span4Mux_h I__2399 (
            .O(N__13221),
            .I(N__13211));
    InMux I__2398 (
            .O(N__13220),
            .I(N__13204));
    InMux I__2397 (
            .O(N__13219),
            .I(N__13204));
    InMux I__2396 (
            .O(N__13216),
            .I(N__13204));
    InMux I__2395 (
            .O(N__13215),
            .I(N__13199));
    InMux I__2394 (
            .O(N__13214),
            .I(N__13199));
    Odrv4 I__2393 (
            .O(N__13211),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2392 (
            .O(N__13204),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2391 (
            .O(N__13199),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    CascadeMux I__2390 (
            .O(N__13192),
            .I(N__13189));
    InMux I__2389 (
            .O(N__13189),
            .I(N__13186));
    LocalMux I__2388 (
            .O(N__13186),
            .I(N__13183));
    Span4Mux_h I__2387 (
            .O(N__13183),
            .I(N__13180));
    Odrv4 I__2386 (
            .O(N__13180),
            .I(\uu2.mem0.w_addr_6 ));
    InMux I__2385 (
            .O(N__13177),
            .I(N__13167));
    InMux I__2384 (
            .O(N__13176),
            .I(N__13164));
    InMux I__2383 (
            .O(N__13175),
            .I(N__13161));
    InMux I__2382 (
            .O(N__13174),
            .I(N__13152));
    InMux I__2381 (
            .O(N__13173),
            .I(N__13152));
    InMux I__2380 (
            .O(N__13172),
            .I(N__13152));
    InMux I__2379 (
            .O(N__13171),
            .I(N__13147));
    InMux I__2378 (
            .O(N__13170),
            .I(N__13147));
    LocalMux I__2377 (
            .O(N__13167),
            .I(N__13142));
    LocalMux I__2376 (
            .O(N__13164),
            .I(N__13142));
    LocalMux I__2375 (
            .O(N__13161),
            .I(N__13139));
    InMux I__2374 (
            .O(N__13160),
            .I(N__13134));
    InMux I__2373 (
            .O(N__13159),
            .I(N__13134));
    LocalMux I__2372 (
            .O(N__13152),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2371 (
            .O(N__13147),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2370 (
            .O(N__13142),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2369 (
            .O(N__13139),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2368 (
            .O(N__13134),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__2367 (
            .O(N__13123),
            .I(N__13120));
    InMux I__2366 (
            .O(N__13120),
            .I(N__13117));
    LocalMux I__2365 (
            .O(N__13117),
            .I(N__13114));
    Span4Mux_h I__2364 (
            .O(N__13114),
            .I(N__13111));
    Odrv4 I__2363 (
            .O(N__13111),
            .I(\uu2.mem0.w_addr_4 ));
    InMux I__2362 (
            .O(N__13108),
            .I(N__13105));
    LocalMux I__2361 (
            .O(N__13105),
            .I(N__13096));
    InMux I__2360 (
            .O(N__13104),
            .I(N__13091));
    InMux I__2359 (
            .O(N__13103),
            .I(N__13091));
    InMux I__2358 (
            .O(N__13102),
            .I(N__13082));
    InMux I__2357 (
            .O(N__13101),
            .I(N__13082));
    InMux I__2356 (
            .O(N__13100),
            .I(N__13082));
    InMux I__2355 (
            .O(N__13099),
            .I(N__13082));
    Odrv4 I__2354 (
            .O(N__13096),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2353 (
            .O(N__13091),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2352 (
            .O(N__13082),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    CascadeMux I__2351 (
            .O(N__13075),
            .I(N__13072));
    InMux I__2350 (
            .O(N__13072),
            .I(N__13069));
    LocalMux I__2349 (
            .O(N__13069),
            .I(N__13066));
    Odrv12 I__2348 (
            .O(N__13066),
            .I(\uu2.mem0.w_addr_5 ));
    CascadeMux I__2347 (
            .O(N__13063),
            .I(N__13060));
    InMux I__2346 (
            .O(N__13060),
            .I(N__13057));
    LocalMux I__2345 (
            .O(N__13057),
            .I(N__13054));
    Odrv12 I__2344 (
            .O(N__13054),
            .I(\uu2.mem0.w_addr_7 ));
    CascadeMux I__2343 (
            .O(N__13051),
            .I(\Lab_UT.dictrl.g0_3_3_cascade_ ));
    InMux I__2342 (
            .O(N__13048),
            .I(N__13045));
    LocalMux I__2341 (
            .O(N__13045),
            .I(N__13042));
    Odrv12 I__2340 (
            .O(N__13042),
            .I(\Lab_UT.dictrl.N_72_mux_0 ));
    InMux I__2339 (
            .O(N__13039),
            .I(N__13035));
    InMux I__2338 (
            .O(N__13038),
            .I(N__13032));
    LocalMux I__2337 (
            .O(N__13035),
            .I(N__13029));
    LocalMux I__2336 (
            .O(N__13032),
            .I(N__13025));
    Span4Mux_h I__2335 (
            .O(N__13029),
            .I(N__13019));
    InMux I__2334 (
            .O(N__13028),
            .I(N__13016));
    Span4Mux_h I__2333 (
            .O(N__13025),
            .I(N__13013));
    InMux I__2332 (
            .O(N__13024),
            .I(N__13008));
    InMux I__2331 (
            .O(N__13023),
            .I(N__13008));
    InMux I__2330 (
            .O(N__13022),
            .I(N__13005));
    Odrv4 I__2329 (
            .O(N__13019),
            .I(bu_rx_data_fast_2));
    LocalMux I__2328 (
            .O(N__13016),
            .I(bu_rx_data_fast_2));
    Odrv4 I__2327 (
            .O(N__13013),
            .I(bu_rx_data_fast_2));
    LocalMux I__2326 (
            .O(N__13008),
            .I(bu_rx_data_fast_2));
    LocalMux I__2325 (
            .O(N__13005),
            .I(bu_rx_data_fast_2));
    InMux I__2324 (
            .O(N__12994),
            .I(N__12987));
    InMux I__2323 (
            .O(N__12993),
            .I(N__12984));
    InMux I__2322 (
            .O(N__12992),
            .I(N__12981));
    InMux I__2321 (
            .O(N__12991),
            .I(N__12978));
    InMux I__2320 (
            .O(N__12990),
            .I(N__12975));
    LocalMux I__2319 (
            .O(N__12987),
            .I(bu_rx_data_fast_1));
    LocalMux I__2318 (
            .O(N__12984),
            .I(bu_rx_data_fast_1));
    LocalMux I__2317 (
            .O(N__12981),
            .I(bu_rx_data_fast_1));
    LocalMux I__2316 (
            .O(N__12978),
            .I(bu_rx_data_fast_1));
    LocalMux I__2315 (
            .O(N__12975),
            .I(bu_rx_data_fast_1));
    InMux I__2314 (
            .O(N__12964),
            .I(N__12959));
    InMux I__2313 (
            .O(N__12963),
            .I(N__12953));
    InMux I__2312 (
            .O(N__12962),
            .I(N__12946));
    LocalMux I__2311 (
            .O(N__12959),
            .I(N__12943));
    InMux I__2310 (
            .O(N__12958),
            .I(N__12938));
    InMux I__2309 (
            .O(N__12957),
            .I(N__12938));
    CascadeMux I__2308 (
            .O(N__12956),
            .I(N__12934));
    LocalMux I__2307 (
            .O(N__12953),
            .I(N__12930));
    InMux I__2306 (
            .O(N__12952),
            .I(N__12925));
    InMux I__2305 (
            .O(N__12951),
            .I(N__12925));
    InMux I__2304 (
            .O(N__12950),
            .I(N__12920));
    InMux I__2303 (
            .O(N__12949),
            .I(N__12920));
    LocalMux I__2302 (
            .O(N__12946),
            .I(N__12913));
    Span4Mux_v I__2301 (
            .O(N__12943),
            .I(N__12913));
    LocalMux I__2300 (
            .O(N__12938),
            .I(N__12913));
    InMux I__2299 (
            .O(N__12937),
            .I(N__12906));
    InMux I__2298 (
            .O(N__12934),
            .I(N__12906));
    InMux I__2297 (
            .O(N__12933),
            .I(N__12906));
    Odrv4 I__2296 (
            .O(N__12930),
            .I(bu_rx_data_6));
    LocalMux I__2295 (
            .O(N__12925),
            .I(bu_rx_data_6));
    LocalMux I__2294 (
            .O(N__12920),
            .I(bu_rx_data_6));
    Odrv4 I__2293 (
            .O(N__12913),
            .I(bu_rx_data_6));
    LocalMux I__2292 (
            .O(N__12906),
            .I(bu_rx_data_6));
    InMux I__2291 (
            .O(N__12895),
            .I(N__12890));
    InMux I__2290 (
            .O(N__12894),
            .I(N__12887));
    InMux I__2289 (
            .O(N__12893),
            .I(N__12880));
    LocalMux I__2288 (
            .O(N__12890),
            .I(N__12875));
    LocalMux I__2287 (
            .O(N__12887),
            .I(N__12875));
    InMux I__2286 (
            .O(N__12886),
            .I(N__12872));
    CascadeMux I__2285 (
            .O(N__12885),
            .I(N__12869));
    InMux I__2284 (
            .O(N__12884),
            .I(N__12861));
    InMux I__2283 (
            .O(N__12883),
            .I(N__12858));
    LocalMux I__2282 (
            .O(N__12880),
            .I(N__12851));
    Span4Mux_v I__2281 (
            .O(N__12875),
            .I(N__12851));
    LocalMux I__2280 (
            .O(N__12872),
            .I(N__12851));
    InMux I__2279 (
            .O(N__12869),
            .I(N__12844));
    InMux I__2278 (
            .O(N__12868),
            .I(N__12844));
    InMux I__2277 (
            .O(N__12867),
            .I(N__12844));
    InMux I__2276 (
            .O(N__12866),
            .I(N__12837));
    InMux I__2275 (
            .O(N__12865),
            .I(N__12837));
    InMux I__2274 (
            .O(N__12864),
            .I(N__12837));
    LocalMux I__2273 (
            .O(N__12861),
            .I(bu_rx_data_5));
    LocalMux I__2272 (
            .O(N__12858),
            .I(bu_rx_data_5));
    Odrv4 I__2271 (
            .O(N__12851),
            .I(bu_rx_data_5));
    LocalMux I__2270 (
            .O(N__12844),
            .I(bu_rx_data_5));
    LocalMux I__2269 (
            .O(N__12837),
            .I(bu_rx_data_5));
    InMux I__2268 (
            .O(N__12826),
            .I(N__12822));
    InMux I__2267 (
            .O(N__12825),
            .I(N__12819));
    LocalMux I__2266 (
            .O(N__12822),
            .I(N__12816));
    LocalMux I__2265 (
            .O(N__12819),
            .I(bu_rx_data_fast_6));
    Odrv4 I__2264 (
            .O(N__12816),
            .I(bu_rx_data_fast_6));
    CascadeMux I__2263 (
            .O(N__12811),
            .I(N__12805));
    InMux I__2262 (
            .O(N__12810),
            .I(N__12797));
    InMux I__2261 (
            .O(N__12809),
            .I(N__12797));
    InMux I__2260 (
            .O(N__12808),
            .I(N__12797));
    InMux I__2259 (
            .O(N__12805),
            .I(N__12791));
    InMux I__2258 (
            .O(N__12804),
            .I(N__12791));
    LocalMux I__2257 (
            .O(N__12797),
            .I(N__12788));
    InMux I__2256 (
            .O(N__12796),
            .I(N__12785));
    LocalMux I__2255 (
            .O(N__12791),
            .I(N__12780));
    Span12Mux_v I__2254 (
            .O(N__12788),
            .I(N__12780));
    LocalMux I__2253 (
            .O(N__12785),
            .I(\uu2.N_40 ));
    Odrv12 I__2252 (
            .O(N__12780),
            .I(\uu2.N_40 ));
    CascadeMux I__2251 (
            .O(N__12775),
            .I(\Lab_UT.i8_mux_0_cascade_ ));
    InMux I__2250 (
            .O(N__12772),
            .I(N__12769));
    LocalMux I__2249 (
            .O(N__12769),
            .I(N__12766));
    Odrv4 I__2248 (
            .O(N__12766),
            .I(\Lab_UT.didp.g0_0_2Z0Z_1 ));
    InMux I__2247 (
            .O(N__12763),
            .I(N__12760));
    LocalMux I__2246 (
            .O(N__12760),
            .I(\Lab_UT.dictrl.g0_0_sn ));
    CascadeMux I__2245 (
            .O(N__12757),
            .I(\Lab_UT.dictrl.g1_1_0_1_cascade_ ));
    InMux I__2244 (
            .O(N__12754),
            .I(N__12751));
    LocalMux I__2243 (
            .O(N__12751),
            .I(\Lab_UT.g1 ));
    InMux I__2242 (
            .O(N__12748),
            .I(N__12745));
    LocalMux I__2241 (
            .O(N__12745),
            .I(\Lab_UT.dictrl.g0_0_rn_0 ));
    CascadeMux I__2240 (
            .O(N__12742),
            .I(N__12737));
    InMux I__2239 (
            .O(N__12741),
            .I(N__12734));
    InMux I__2238 (
            .O(N__12740),
            .I(N__12729));
    InMux I__2237 (
            .O(N__12737),
            .I(N__12729));
    LocalMux I__2236 (
            .O(N__12734),
            .I(\Lab_UT.dictrl.m22Z0Z_1 ));
    LocalMux I__2235 (
            .O(N__12729),
            .I(\Lab_UT.dictrl.m22Z0Z_1 ));
    InMux I__2234 (
            .O(N__12724),
            .I(N__12719));
    IoInMux I__2233 (
            .O(N__12723),
            .I(N__12716));
    InMux I__2232 (
            .O(N__12722),
            .I(N__12712));
    LocalMux I__2231 (
            .O(N__12719),
            .I(N__12709));
    LocalMux I__2230 (
            .O(N__12716),
            .I(N__12706));
    InMux I__2229 (
            .O(N__12715),
            .I(N__12703));
    LocalMux I__2228 (
            .O(N__12712),
            .I(N__12700));
    Span4Mux_h I__2227 (
            .O(N__12709),
            .I(N__12697));
    IoSpan4Mux I__2226 (
            .O(N__12706),
            .I(N__12694));
    LocalMux I__2225 (
            .O(N__12703),
            .I(N__12691));
    Span4Mux_h I__2224 (
            .O(N__12700),
            .I(N__12688));
    Span4Mux_h I__2223 (
            .O(N__12697),
            .I(N__12683));
    Span4Mux_s1_h I__2222 (
            .O(N__12694),
            .I(N__12683));
    Odrv12 I__2221 (
            .O(N__12691),
            .I(rst));
    Odrv4 I__2220 (
            .O(N__12688),
            .I(rst));
    Odrv4 I__2219 (
            .O(N__12683),
            .I(rst));
    CascadeMux I__2218 (
            .O(N__12676),
            .I(\Lab_UT.dictrl.g1_1_0_0_cascade_ ));
    InMux I__2217 (
            .O(N__12673),
            .I(N__12670));
    LocalMux I__2216 (
            .O(N__12670),
            .I(\Lab_UT.dictrl.g1_1_0 ));
    InMux I__2215 (
            .O(N__12667),
            .I(N__12664));
    LocalMux I__2214 (
            .O(N__12664),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1 ));
    InMux I__2213 (
            .O(N__12661),
            .I(N__12658));
    LocalMux I__2212 (
            .O(N__12658),
            .I(\Lab_UT.dictrl.N_3 ));
    CascadeMux I__2211 (
            .O(N__12655),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ));
    InMux I__2210 (
            .O(N__12652),
            .I(N__12649));
    LocalMux I__2209 (
            .O(N__12649),
            .I(\Lab_UT.dictrl.m37_N_2LZ0Z1 ));
    InMux I__2208 (
            .O(N__12646),
            .I(N__12643));
    LocalMux I__2207 (
            .O(N__12643),
            .I(\Lab_UT.dictrl.N_72_mux_1 ));
    CascadeMux I__2206 (
            .O(N__12640),
            .I(\Lab_UT.dictrl.G_25_i_1_cascade_ ));
    InMux I__2205 (
            .O(N__12637),
            .I(N__12634));
    LocalMux I__2204 (
            .O(N__12634),
            .I(\Lab_UT.dictrl.G_25_i_0 ));
    InMux I__2203 (
            .O(N__12631),
            .I(N__12628));
    LocalMux I__2202 (
            .O(N__12628),
            .I(\Lab_UT.dictrl.G_25_i_a5_1_0 ));
    CascadeMux I__2201 (
            .O(N__12625),
            .I(\Lab_UT.dictrl.N_18_0_0_cascade_ ));
    InMux I__2200 (
            .O(N__12622),
            .I(N__12619));
    LocalMux I__2199 (
            .O(N__12619),
            .I(\Lab_UT.dictrl.g0_6_3_0 ));
    CascadeMux I__2198 (
            .O(N__12616),
            .I(N__12613));
    InMux I__2197 (
            .O(N__12613),
            .I(N__12610));
    LocalMux I__2196 (
            .O(N__12610),
            .I(N__12607));
    Odrv12 I__2195 (
            .O(N__12607),
            .I(\Lab_UT.dictrl.g2Z0Z_0 ));
    CascadeMux I__2194 (
            .O(N__12604),
            .I(N__12600));
    InMux I__2193 (
            .O(N__12603),
            .I(N__12596));
    InMux I__2192 (
            .O(N__12600),
            .I(N__12593));
    InMux I__2191 (
            .O(N__12599),
            .I(N__12590));
    LocalMux I__2190 (
            .O(N__12596),
            .I(\Lab_UT.dispString.N_145 ));
    LocalMux I__2189 (
            .O(N__12593),
            .I(\Lab_UT.dispString.N_145 ));
    LocalMux I__2188 (
            .O(N__12590),
            .I(\Lab_UT.dispString.N_145 ));
    CascadeMux I__2187 (
            .O(N__12583),
            .I(\Lab_UT.dispString.N_118_cascade_ ));
    InMux I__2186 (
            .O(N__12580),
            .I(N__12577));
    LocalMux I__2185 (
            .O(N__12577),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_1 ));
    CEMux I__2184 (
            .O(N__12574),
            .I(N__12571));
    LocalMux I__2183 (
            .O(N__12571),
            .I(N__12568));
    Span4Mux_v I__2182 (
            .O(N__12568),
            .I(N__12564));
    CEMux I__2181 (
            .O(N__12567),
            .I(N__12561));
    Span4Mux_v I__2180 (
            .O(N__12564),
            .I(N__12556));
    LocalMux I__2179 (
            .O(N__12561),
            .I(N__12556));
    Span4Mux_v I__2178 (
            .O(N__12556),
            .I(N__12553));
    Sp12to4 I__2177 (
            .O(N__12553),
            .I(N__12550));
    Odrv12 I__2176 (
            .O(N__12550),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    InMux I__2175 (
            .O(N__12547),
            .I(N__12544));
    LocalMux I__2174 (
            .O(N__12544),
            .I(N__12541));
    Span4Mux_v I__2173 (
            .O(N__12541),
            .I(N__12538));
    Odrv4 I__2172 (
            .O(N__12538),
            .I(\Lab_UT.dictrl.G_25_i_o3_4 ));
    InMux I__2171 (
            .O(N__12535),
            .I(N__12532));
    LocalMux I__2170 (
            .O(N__12532),
            .I(\Lab_UT.dictrl.G_25_i_o3_5 ));
    CascadeMux I__2169 (
            .O(N__12529),
            .I(\Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ));
    CascadeMux I__2168 (
            .O(N__12526),
            .I(\Lab_UT.dictrl.N_11_cascade_ ));
    CascadeMux I__2167 (
            .O(N__12523),
            .I(N__12520));
    InMux I__2166 (
            .O(N__12520),
            .I(N__12512));
    InMux I__2165 (
            .O(N__12519),
            .I(N__12512));
    InMux I__2164 (
            .O(N__12518),
            .I(N__12507));
    InMux I__2163 (
            .O(N__12517),
            .I(N__12507));
    LocalMux I__2162 (
            .O(N__12512),
            .I(N__12504));
    LocalMux I__2161 (
            .O(N__12507),
            .I(N__12501));
    Span4Mux_h I__2160 (
            .O(N__12504),
            .I(N__12496));
    Span4Mux_v I__2159 (
            .O(N__12501),
            .I(N__12496));
    Odrv4 I__2158 (
            .O(N__12496),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    CascadeMux I__2157 (
            .O(N__12493),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_ ));
    InMux I__2156 (
            .O(N__12490),
            .I(N__12486));
    InMux I__2155 (
            .O(N__12489),
            .I(N__12483));
    LocalMux I__2154 (
            .O(N__12486),
            .I(N__12479));
    LocalMux I__2153 (
            .O(N__12483),
            .I(N__12476));
    InMux I__2152 (
            .O(N__12482),
            .I(N__12473));
    Span4Mux_h I__2151 (
            .O(N__12479),
            .I(N__12470));
    Span4Mux_v I__2150 (
            .O(N__12476),
            .I(N__12465));
    LocalMux I__2149 (
            .O(N__12473),
            .I(N__12465));
    Odrv4 I__2148 (
            .O(N__12470),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv4 I__2147 (
            .O(N__12465),
            .I(\Lab_UT.di_AStens_3 ));
    CascadeMux I__2146 (
            .O(N__12460),
            .I(N__12453));
    InMux I__2145 (
            .O(N__12459),
            .I(N__12450));
    InMux I__2144 (
            .O(N__12458),
            .I(N__12447));
    InMux I__2143 (
            .O(N__12457),
            .I(N__12442));
    InMux I__2142 (
            .O(N__12456),
            .I(N__12442));
    InMux I__2141 (
            .O(N__12453),
            .I(N__12439));
    LocalMux I__2140 (
            .O(N__12450),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2139 (
            .O(N__12447),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2138 (
            .O(N__12442),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2137 (
            .O(N__12439),
            .I(\Lab_UT.di_Stens_3 ));
    InMux I__2136 (
            .O(N__12430),
            .I(N__12427));
    LocalMux I__2135 (
            .O(N__12427),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ));
    CascadeMux I__2134 (
            .O(N__12424),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_ ));
    InMux I__2133 (
            .O(N__12421),
            .I(N__12418));
    LocalMux I__2132 (
            .O(N__12418),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0 ));
    InMux I__2131 (
            .O(N__12415),
            .I(N__12412));
    LocalMux I__2130 (
            .O(N__12412),
            .I(N__12409));
    Odrv4 I__2129 (
            .O(N__12409),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ));
    CascadeMux I__2128 (
            .O(N__12406),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ));
    InMux I__2127 (
            .O(N__12403),
            .I(N__12400));
    LocalMux I__2126 (
            .O(N__12400),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ));
    InMux I__2125 (
            .O(N__12397),
            .I(N__12391));
    InMux I__2124 (
            .O(N__12396),
            .I(N__12384));
    InMux I__2123 (
            .O(N__12395),
            .I(N__12384));
    InMux I__2122 (
            .O(N__12394),
            .I(N__12384));
    LocalMux I__2121 (
            .O(N__12391),
            .I(N__12379));
    LocalMux I__2120 (
            .O(N__12384),
            .I(N__12379));
    Span4Mux_h I__2119 (
            .O(N__12379),
            .I(N__12376));
    Odrv4 I__2118 (
            .O(N__12376),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ));
    InMux I__2117 (
            .O(N__12373),
            .I(N__12370));
    LocalMux I__2116 (
            .O(N__12370),
            .I(N__12365));
    InMux I__2115 (
            .O(N__12369),
            .I(N__12362));
    InMux I__2114 (
            .O(N__12368),
            .I(N__12359));
    Span4Mux_v I__2113 (
            .O(N__12365),
            .I(N__12354));
    LocalMux I__2112 (
            .O(N__12362),
            .I(N__12354));
    LocalMux I__2111 (
            .O(N__12359),
            .I(\Lab_UT.di_AStens_0 ));
    Odrv4 I__2110 (
            .O(N__12354),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__2109 (
            .O(N__12349),
            .I(N__12346));
    LocalMux I__2108 (
            .O(N__12346),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ));
    CascadeMux I__2107 (
            .O(N__12343),
            .I(\Lab_UT.didp.countrce4.q_5_0_cascade_ ));
    InMux I__2106 (
            .O(N__12340),
            .I(N__12336));
    CascadeMux I__2105 (
            .O(N__12339),
            .I(N__12333));
    LocalMux I__2104 (
            .O(N__12336),
            .I(N__12330));
    InMux I__2103 (
            .O(N__12333),
            .I(N__12327));
    Span4Mux_v I__2102 (
            .O(N__12330),
            .I(N__12324));
    LocalMux I__2101 (
            .O(N__12327),
            .I(N__12321));
    Odrv4 I__2100 (
            .O(N__12324),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv12 I__2099 (
            .O(N__12321),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    CEMux I__2098 (
            .O(N__12316),
            .I(N__12313));
    LocalMux I__2097 (
            .O(N__12313),
            .I(N__12310));
    Span4Mux_v I__2096 (
            .O(N__12310),
            .I(N__12307));
    Span4Mux_h I__2095 (
            .O(N__12307),
            .I(N__12304));
    Odrv4 I__2094 (
            .O(N__12304),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    CascadeMux I__2093 (
            .O(N__12301),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_ ));
    InMux I__2092 (
            .O(N__12298),
            .I(N__12295));
    LocalMux I__2091 (
            .O(N__12295),
            .I(N__12292));
    Odrv4 I__2090 (
            .O(N__12292),
            .I(\Lab_UT.didp.countrce2.N_96 ));
    CascadeMux I__2089 (
            .O(N__12289),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_ ));
    InMux I__2088 (
            .O(N__12286),
            .I(N__12282));
    InMux I__2087 (
            .O(N__12285),
            .I(N__12278));
    LocalMux I__2086 (
            .O(N__12282),
            .I(N__12275));
    InMux I__2085 (
            .O(N__12281),
            .I(N__12272));
    LocalMux I__2084 (
            .O(N__12278),
            .I(N__12269));
    Span4Mux_v I__2083 (
            .O(N__12275),
            .I(N__12266));
    LocalMux I__2082 (
            .O(N__12272),
            .I(N__12263));
    Odrv4 I__2081 (
            .O(N__12269),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__2080 (
            .O(N__12266),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__2079 (
            .O(N__12263),
            .I(\Lab_UT.di_AStens_2 ));
    CascadeMux I__2078 (
            .O(N__12256),
            .I(N__12249));
    CascadeMux I__2077 (
            .O(N__12255),
            .I(N__12245));
    InMux I__2076 (
            .O(N__12254),
            .I(N__12234));
    InMux I__2075 (
            .O(N__12253),
            .I(N__12234));
    InMux I__2074 (
            .O(N__12252),
            .I(N__12234));
    InMux I__2073 (
            .O(N__12249),
            .I(N__12234));
    InMux I__2072 (
            .O(N__12248),
            .I(N__12234));
    InMux I__2071 (
            .O(N__12245),
            .I(N__12231));
    LocalMux I__2070 (
            .O(N__12234),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__2069 (
            .O(N__12231),
            .I(\Lab_UT.di_Stens_2 ));
    CascadeMux I__2068 (
            .O(N__12226),
            .I(N__12221));
    InMux I__2067 (
            .O(N__12225),
            .I(N__12218));
    InMux I__2066 (
            .O(N__12224),
            .I(N__12215));
    InMux I__2065 (
            .O(N__12221),
            .I(N__12212));
    LocalMux I__2064 (
            .O(N__12218),
            .I(N__12209));
    LocalMux I__2063 (
            .O(N__12215),
            .I(N__12206));
    LocalMux I__2062 (
            .O(N__12212),
            .I(N__12203));
    Span4Mux_h I__2061 (
            .O(N__12209),
            .I(N__12200));
    Span4Mux_h I__2060 (
            .O(N__12206),
            .I(N__12197));
    Odrv12 I__2059 (
            .O(N__12203),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__2058 (
            .O(N__12200),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__2057 (
            .O(N__12197),
            .I(\Lab_UT.di_AMones_0 ));
    InMux I__2056 (
            .O(N__12190),
            .I(N__12187));
    LocalMux I__2055 (
            .O(N__12187),
            .I(N__12184));
    Span4Mux_h I__2054 (
            .O(N__12184),
            .I(N__12181));
    Odrv4 I__2053 (
            .O(N__12181),
            .I(\uu2.bitmapZ0Z_180 ));
    InMux I__2052 (
            .O(N__12178),
            .I(N__12175));
    LocalMux I__2051 (
            .O(N__12175),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__2050 (
            .O(N__12172),
            .I(N__12169));
    LocalMux I__2049 (
            .O(N__12169),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__2048 (
            .O(N__12166),
            .I(N__12163));
    LocalMux I__2047 (
            .O(N__12163),
            .I(N__12160));
    Span4Mux_h I__2046 (
            .O(N__12160),
            .I(N__12157));
    Odrv4 I__2045 (
            .O(N__12157),
            .I(\uu2.N_149 ));
    InMux I__2044 (
            .O(N__12154),
            .I(N__12151));
    LocalMux I__2043 (
            .O(N__12151),
            .I(\uu2.bitmapZ0Z_84 ));
    CascadeMux I__2042 (
            .O(N__12148),
            .I(N__12145));
    InMux I__2041 (
            .O(N__12145),
            .I(N__12142));
    LocalMux I__2040 (
            .O(N__12142),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__2039 (
            .O(N__12139),
            .I(N__12136));
    LocalMux I__2038 (
            .O(N__12136),
            .I(\uu2.N_25 ));
    CascadeMux I__2037 (
            .O(N__12133),
            .I(N__12130));
    InMux I__2036 (
            .O(N__12130),
            .I(N__12124));
    InMux I__2035 (
            .O(N__12129),
            .I(N__12124));
    LocalMux I__2034 (
            .O(N__12124),
            .I(N__12118));
    InMux I__2033 (
            .O(N__12123),
            .I(N__12111));
    InMux I__2032 (
            .O(N__12122),
            .I(N__12111));
    InMux I__2031 (
            .O(N__12121),
            .I(N__12111));
    Odrv12 I__2030 (
            .O(N__12118),
            .I(\Lab_UT.didp.un24_ce_3 ));
    LocalMux I__2029 (
            .O(N__12111),
            .I(\Lab_UT.didp.un24_ce_3 ));
    CascadeMux I__2028 (
            .O(N__12106),
            .I(N__12098));
    InMux I__2027 (
            .O(N__12105),
            .I(N__12094));
    InMux I__2026 (
            .O(N__12104),
            .I(N__12091));
    InMux I__2025 (
            .O(N__12103),
            .I(N__12080));
    InMux I__2024 (
            .O(N__12102),
            .I(N__12080));
    InMux I__2023 (
            .O(N__12101),
            .I(N__12080));
    InMux I__2022 (
            .O(N__12098),
            .I(N__12080));
    InMux I__2021 (
            .O(N__12097),
            .I(N__12080));
    LocalMux I__2020 (
            .O(N__12094),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2019 (
            .O(N__12091),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2018 (
            .O(N__12080),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    InMux I__2017 (
            .O(N__12073),
            .I(N__12070));
    LocalMux I__2016 (
            .O(N__12070),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__2015 (
            .O(N__12067),
            .I(N__12064));
    InMux I__2014 (
            .O(N__12064),
            .I(N__12061));
    LocalMux I__2013 (
            .O(N__12061),
            .I(N__12058));
    Odrv4 I__2012 (
            .O(N__12058),
            .I(\uu2.bitmapZ0Z_221 ));
    InMux I__2011 (
            .O(N__12055),
            .I(N__12052));
    LocalMux I__2010 (
            .O(N__12052),
            .I(\uu2.bitmapZ0Z_75 ));
    CascadeMux I__2009 (
            .O(N__12049),
            .I(N__12046));
    InMux I__2008 (
            .O(N__12046),
            .I(N__12043));
    LocalMux I__2007 (
            .O(N__12043),
            .I(\uu2.bitmapZ0Z_203 ));
    CascadeMux I__2006 (
            .O(N__12040),
            .I(\uu2.N_24_cascade_ ));
    InMux I__2005 (
            .O(N__12037),
            .I(N__12031));
    InMux I__2004 (
            .O(N__12036),
            .I(N__12031));
    LocalMux I__2003 (
            .O(N__12031),
            .I(\uu2.N_31_i ));
    InMux I__2002 (
            .O(N__12028),
            .I(N__12025));
    LocalMux I__2001 (
            .O(N__12025),
            .I(\uu2.N_166 ));
    CascadeMux I__2000 (
            .O(N__12022),
            .I(\uu2.bitmap_pmux_27_ns_1_cascade_ ));
    InMux I__1999 (
            .O(N__12019),
            .I(N__12016));
    LocalMux I__1998 (
            .O(N__12016),
            .I(\uu2.N_26 ));
    InMux I__1997 (
            .O(N__12013),
            .I(N__12010));
    LocalMux I__1996 (
            .O(N__12010),
            .I(N__12007));
    Span4Mux_s2_v I__1995 (
            .O(N__12007),
            .I(N__12004));
    Odrv4 I__1994 (
            .O(N__12004),
            .I(\uu2.N_404 ));
    InMux I__1993 (
            .O(N__12001),
            .I(N__11998));
    LocalMux I__1992 (
            .O(N__11998),
            .I(N__11995));
    Span4Mux_h I__1991 (
            .O(N__11995),
            .I(N__11992));
    Odrv4 I__1990 (
            .O(N__11992),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    InMux I__1989 (
            .O(N__11989),
            .I(N__11983));
    InMux I__1988 (
            .O(N__11988),
            .I(N__11978));
    InMux I__1987 (
            .O(N__11987),
            .I(N__11978));
    InMux I__1986 (
            .O(N__11986),
            .I(N__11975));
    LocalMux I__1985 (
            .O(N__11983),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__1984 (
            .O(N__11978),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__1983 (
            .O(N__11975),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__1982 (
            .O(N__11968),
            .I(N__11965));
    LocalMux I__1981 (
            .O(N__11965),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    CascadeMux I__1980 (
            .O(N__11962),
            .I(\uu2.N_14_cascade_ ));
    InMux I__1979 (
            .O(N__11959),
            .I(N__11956));
    LocalMux I__1978 (
            .O(N__11956),
            .I(\uu2.bitmap_pmux_sn_N_54_mux ));
    InMux I__1977 (
            .O(N__11953),
            .I(N__11950));
    LocalMux I__1976 (
            .O(N__11950),
            .I(\uu2.bitmap_RNI2Q8F1Z0Z_111 ));
    InMux I__1975 (
            .O(N__11947),
            .I(N__11940));
    InMux I__1974 (
            .O(N__11946),
            .I(N__11933));
    InMux I__1973 (
            .O(N__11945),
            .I(N__11933));
    InMux I__1972 (
            .O(N__11944),
            .I(N__11933));
    InMux I__1971 (
            .O(N__11943),
            .I(N__11930));
    LocalMux I__1970 (
            .O(N__11940),
            .I(N__11927));
    LocalMux I__1969 (
            .O(N__11933),
            .I(N__11924));
    LocalMux I__1968 (
            .O(N__11930),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__1967 (
            .O(N__11927),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__1966 (
            .O(N__11924),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__1965 (
            .O(N__11917),
            .I(N__11914));
    LocalMux I__1964 (
            .O(N__11914),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__1963 (
            .O(N__11911),
            .I(N__11907));
    InMux I__1962 (
            .O(N__11910),
            .I(N__11902));
    InMux I__1961 (
            .O(N__11907),
            .I(N__11902));
    LocalMux I__1960 (
            .O(N__11902),
            .I(bu_rx_data_fast_5));
    CascadeMux I__1959 (
            .O(N__11899),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ));
    CascadeMux I__1958 (
            .O(N__11896),
            .I(N__11890));
    CascadeMux I__1957 (
            .O(N__11895),
            .I(N__11887));
    CascadeMux I__1956 (
            .O(N__11894),
            .I(N__11883));
    CascadeMux I__1955 (
            .O(N__11893),
            .I(N__11878));
    InMux I__1954 (
            .O(N__11890),
            .I(N__11875));
    InMux I__1953 (
            .O(N__11887),
            .I(N__11862));
    InMux I__1952 (
            .O(N__11886),
            .I(N__11862));
    InMux I__1951 (
            .O(N__11883),
            .I(N__11862));
    InMux I__1950 (
            .O(N__11882),
            .I(N__11862));
    InMux I__1949 (
            .O(N__11881),
            .I(N__11862));
    InMux I__1948 (
            .O(N__11878),
            .I(N__11862));
    LocalMux I__1947 (
            .O(N__11875),
            .I(N__11859));
    LocalMux I__1946 (
            .O(N__11862),
            .I(N__11856));
    Span4Mux_h I__1945 (
            .O(N__11859),
            .I(N__11851));
    Span4Mux_s0_v I__1944 (
            .O(N__11856),
            .I(N__11851));
    Odrv4 I__1943 (
            .O(N__11851),
            .I(\uu2.N_37 ));
    InMux I__1942 (
            .O(N__11848),
            .I(N__11845));
    LocalMux I__1941 (
            .O(N__11845),
            .I(N__11842));
    Odrv4 I__1940 (
            .O(N__11842),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    CascadeMux I__1939 (
            .O(N__11839),
            .I(\resetGen.escKeyZ0Z_4_cascade_ ));
    InMux I__1938 (
            .O(N__11836),
            .I(N__11821));
    InMux I__1937 (
            .O(N__11835),
            .I(N__11821));
    InMux I__1936 (
            .O(N__11834),
            .I(N__11821));
    InMux I__1935 (
            .O(N__11833),
            .I(N__11821));
    InMux I__1934 (
            .O(N__11832),
            .I(N__11821));
    LocalMux I__1933 (
            .O(N__11821),
            .I(N__11818));
    Span4Mux_h I__1932 (
            .O(N__11818),
            .I(N__11815));
    Odrv4 I__1931 (
            .O(N__11815),
            .I(\resetGen.escKeyZ0 ));
    InMux I__1930 (
            .O(N__11812),
            .I(N__11809));
    LocalMux I__1929 (
            .O(N__11809),
            .I(\resetGen.escKeyZ0Z_5 ));
    InMux I__1928 (
            .O(N__11806),
            .I(N__11803));
    LocalMux I__1927 (
            .O(N__11803),
            .I(\Lab_UT.dictrl.g1_0Z0Z_5 ));
    InMux I__1926 (
            .O(N__11800),
            .I(N__11797));
    LocalMux I__1925 (
            .O(N__11797),
            .I(N__11794));
    Odrv4 I__1924 (
            .O(N__11794),
            .I(\Lab_UT.dictrl.g1_4_0 ));
    CascadeMux I__1923 (
            .O(N__11791),
            .I(\Lab_UT.dictrl.g1_5_0_cascade_ ));
    CascadeMux I__1922 (
            .O(N__11788),
            .I(\Lab_UT.dictrl.G_25_i_o3_3_cascade_ ));
    InMux I__1921 (
            .O(N__11785),
            .I(N__11782));
    LocalMux I__1920 (
            .O(N__11782),
            .I(\Lab_UT.dictrl.g0_5_3_0 ));
    CascadeMux I__1919 (
            .O(N__11779),
            .I(\Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ));
    InMux I__1918 (
            .O(N__11776),
            .I(N__11771));
    InMux I__1917 (
            .O(N__11775),
            .I(N__11768));
    InMux I__1916 (
            .O(N__11774),
            .I(N__11765));
    LocalMux I__1915 (
            .O(N__11771),
            .I(\Lab_UT.dispString.N_144 ));
    LocalMux I__1914 (
            .O(N__11768),
            .I(\Lab_UT.dispString.N_144 ));
    LocalMux I__1913 (
            .O(N__11765),
            .I(\Lab_UT.dispString.N_144 ));
    InMux I__1912 (
            .O(N__11758),
            .I(N__11755));
    LocalMux I__1911 (
            .O(N__11755),
            .I(\Lab_UT.dispString.N_124 ));
    CascadeMux I__1910 (
            .O(N__11752),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_ ));
    InMux I__1909 (
            .O(N__11749),
            .I(N__11743));
    InMux I__1908 (
            .O(N__11748),
            .I(N__11740));
    InMux I__1907 (
            .O(N__11747),
            .I(N__11737));
    InMux I__1906 (
            .O(N__11746),
            .I(N__11734));
    LocalMux I__1905 (
            .O(N__11743),
            .I(N__11731));
    LocalMux I__1904 (
            .O(N__11740),
            .I(\Lab_UT.dispString.N_95 ));
    LocalMux I__1903 (
            .O(N__11737),
            .I(\Lab_UT.dispString.N_95 ));
    LocalMux I__1902 (
            .O(N__11734),
            .I(\Lab_UT.dispString.N_95 ));
    Odrv4 I__1901 (
            .O(N__11731),
            .I(\Lab_UT.dispString.N_95 ));
    InMux I__1900 (
            .O(N__11722),
            .I(N__11719));
    LocalMux I__1899 (
            .O(N__11719),
            .I(\Lab_UT.dispString.N_102 ));
    CascadeMux I__1898 (
            .O(N__11716),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ));
    InMux I__1897 (
            .O(N__11713),
            .I(N__11710));
    LocalMux I__1896 (
            .O(N__11710),
            .I(N__11707));
    Span4Mux_h I__1895 (
            .O(N__11707),
            .I(N__11704));
    Span4Mux_v I__1894 (
            .O(N__11704),
            .I(N__11699));
    InMux I__1893 (
            .O(N__11703),
            .I(N__11694));
    InMux I__1892 (
            .O(N__11702),
            .I(N__11694));
    Odrv4 I__1891 (
            .O(N__11699),
            .I(L3_tx_data_0));
    LocalMux I__1890 (
            .O(N__11694),
            .I(L3_tx_data_0));
    InMux I__1889 (
            .O(N__11689),
            .I(N__11681));
    InMux I__1888 (
            .O(N__11688),
            .I(N__11681));
    InMux I__1887 (
            .O(N__11687),
            .I(N__11678));
    InMux I__1886 (
            .O(N__11686),
            .I(N__11675));
    LocalMux I__1885 (
            .O(N__11681),
            .I(N__11672));
    LocalMux I__1884 (
            .O(N__11678),
            .I(\Lab_UT.dispString.N_143 ));
    LocalMux I__1883 (
            .O(N__11675),
            .I(\Lab_UT.dispString.N_143 ));
    Odrv4 I__1882 (
            .O(N__11672),
            .I(\Lab_UT.dispString.N_143 ));
    CascadeMux I__1881 (
            .O(N__11665),
            .I(N__11661));
    CascadeMux I__1880 (
            .O(N__11664),
            .I(N__11658));
    InMux I__1879 (
            .O(N__11661),
            .I(N__11650));
    InMux I__1878 (
            .O(N__11658),
            .I(N__11647));
    InMux I__1877 (
            .O(N__11657),
            .I(N__11642));
    InMux I__1876 (
            .O(N__11656),
            .I(N__11642));
    CascadeMux I__1875 (
            .O(N__11655),
            .I(N__11638));
    CascadeMux I__1874 (
            .O(N__11654),
            .I(N__11634));
    CascadeMux I__1873 (
            .O(N__11653),
            .I(N__11631));
    LocalMux I__1872 (
            .O(N__11650),
            .I(N__11626));
    LocalMux I__1871 (
            .O(N__11647),
            .I(N__11626));
    LocalMux I__1870 (
            .O(N__11642),
            .I(N__11623));
    InMux I__1869 (
            .O(N__11641),
            .I(N__11618));
    InMux I__1868 (
            .O(N__11638),
            .I(N__11618));
    InMux I__1867 (
            .O(N__11637),
            .I(N__11611));
    InMux I__1866 (
            .O(N__11634),
            .I(N__11611));
    InMux I__1865 (
            .O(N__11631),
            .I(N__11611));
    Span4Mux_v I__1864 (
            .O(N__11626),
            .I(N__11608));
    Odrv4 I__1863 (
            .O(N__11623),
            .I(oneSecStrb));
    LocalMux I__1862 (
            .O(N__11618),
            .I(oneSecStrb));
    LocalMux I__1861 (
            .O(N__11611),
            .I(oneSecStrb));
    Odrv4 I__1860 (
            .O(N__11608),
            .I(oneSecStrb));
    InMux I__1859 (
            .O(N__11599),
            .I(N__11596));
    LocalMux I__1858 (
            .O(N__11596),
            .I(N__11593));
    Span4Mux_h I__1857 (
            .O(N__11593),
            .I(N__11590));
    Odrv4 I__1856 (
            .O(N__11590),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_1 ));
    CEMux I__1855 (
            .O(N__11587),
            .I(N__11584));
    LocalMux I__1854 (
            .O(N__11584),
            .I(N__11581));
    Span4Mux_h I__1853 (
            .O(N__11581),
            .I(N__11578));
    Odrv4 I__1852 (
            .O(N__11578),
            .I(\Lab_UT.didp.regrce2.LdAStens_0 ));
    InMux I__1851 (
            .O(N__11575),
            .I(N__11568));
    InMux I__1850 (
            .O(N__11574),
            .I(N__11568));
    InMux I__1849 (
            .O(N__11573),
            .I(N__11562));
    LocalMux I__1848 (
            .O(N__11568),
            .I(N__11559));
    InMux I__1847 (
            .O(N__11567),
            .I(N__11552));
    InMux I__1846 (
            .O(N__11566),
            .I(N__11552));
    InMux I__1845 (
            .O(N__11565),
            .I(N__11552));
    LocalMux I__1844 (
            .O(N__11562),
            .I(N__11549));
    Span4Mux_h I__1843 (
            .O(N__11559),
            .I(N__11544));
    LocalMux I__1842 (
            .O(N__11552),
            .I(N__11544));
    Odrv12 I__1841 (
            .O(N__11549),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    Odrv4 I__1840 (
            .O(N__11544),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    CascadeMux I__1839 (
            .O(N__11539),
            .I(\Lab_UT.dispString.N_102_cascade_ ));
    InMux I__1838 (
            .O(N__11536),
            .I(N__11533));
    LocalMux I__1837 (
            .O(N__11533),
            .I(N__11529));
    InMux I__1836 (
            .O(N__11532),
            .I(N__11526));
    Odrv4 I__1835 (
            .O(N__11529),
            .I(G_186));
    LocalMux I__1834 (
            .O(N__11526),
            .I(G_186));
    InMux I__1833 (
            .O(N__11521),
            .I(N__11518));
    LocalMux I__1832 (
            .O(N__11518),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_2 ));
    CascadeMux I__1831 (
            .O(N__11515),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_ ));
    InMux I__1830 (
            .O(N__11512),
            .I(N__11509));
    LocalMux I__1829 (
            .O(N__11509),
            .I(N__11505));
    CascadeMux I__1828 (
            .O(N__11508),
            .I(N__11501));
    Span4Mux_v I__1827 (
            .O(N__11505),
            .I(N__11498));
    InMux I__1826 (
            .O(N__11504),
            .I(N__11493));
    InMux I__1825 (
            .O(N__11501),
            .I(N__11493));
    Odrv4 I__1824 (
            .O(N__11498),
            .I(L3_tx_data_2));
    LocalMux I__1823 (
            .O(N__11493),
            .I(L3_tx_data_2));
    InMux I__1822 (
            .O(N__11488),
            .I(N__11484));
    InMux I__1821 (
            .O(N__11487),
            .I(N__11481));
    LocalMux I__1820 (
            .O(N__11484),
            .I(N__11478));
    LocalMux I__1819 (
            .O(N__11481),
            .I(N__11472));
    Span4Mux_s3_v I__1818 (
            .O(N__11478),
            .I(N__11472));
    InMux I__1817 (
            .O(N__11477),
            .I(N__11469));
    Odrv4 I__1816 (
            .O(N__11472),
            .I(L3_tx_data_rdy));
    LocalMux I__1815 (
            .O(N__11469),
            .I(L3_tx_data_rdy));
    InMux I__1814 (
            .O(N__11464),
            .I(N__11461));
    LocalMux I__1813 (
            .O(N__11461),
            .I(N__11456));
    InMux I__1812 (
            .O(N__11460),
            .I(N__11453));
    InMux I__1811 (
            .O(N__11459),
            .I(N__11450));
    Odrv4 I__1810 (
            .O(N__11456),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    LocalMux I__1809 (
            .O(N__11453),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    LocalMux I__1808 (
            .O(N__11450),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    InMux I__1807 (
            .O(N__11443),
            .I(N__11440));
    LocalMux I__1806 (
            .O(N__11440),
            .I(N__11435));
    InMux I__1805 (
            .O(N__11439),
            .I(N__11432));
    InMux I__1804 (
            .O(N__11438),
            .I(N__11429));
    Odrv4 I__1803 (
            .O(N__11435),
            .I(\uu2.un1_w_user_crZ0Z_3 ));
    LocalMux I__1802 (
            .O(N__11432),
            .I(\uu2.un1_w_user_crZ0Z_3 ));
    LocalMux I__1801 (
            .O(N__11429),
            .I(\uu2.un1_w_user_crZ0Z_3 ));
    InMux I__1800 (
            .O(N__11422),
            .I(N__11419));
    LocalMux I__1799 (
            .O(N__11419),
            .I(N__11416));
    Span4Mux_v I__1798 (
            .O(N__11416),
            .I(N__11404));
    InMux I__1797 (
            .O(N__11415),
            .I(N__11401));
    InMux I__1796 (
            .O(N__11414),
            .I(N__11398));
    InMux I__1795 (
            .O(N__11413),
            .I(N__11395));
    InMux I__1794 (
            .O(N__11412),
            .I(N__11392));
    InMux I__1793 (
            .O(N__11411),
            .I(N__11387));
    InMux I__1792 (
            .O(N__11410),
            .I(N__11387));
    InMux I__1791 (
            .O(N__11409),
            .I(N__11380));
    InMux I__1790 (
            .O(N__11408),
            .I(N__11380));
    InMux I__1789 (
            .O(N__11407),
            .I(N__11380));
    Odrv4 I__1788 (
            .O(N__11404),
            .I(G_179));
    LocalMux I__1787 (
            .O(N__11401),
            .I(G_179));
    LocalMux I__1786 (
            .O(N__11398),
            .I(G_179));
    LocalMux I__1785 (
            .O(N__11395),
            .I(G_179));
    LocalMux I__1784 (
            .O(N__11392),
            .I(G_179));
    LocalMux I__1783 (
            .O(N__11387),
            .I(G_179));
    LocalMux I__1782 (
            .O(N__11380),
            .I(G_179));
    CascadeMux I__1781 (
            .O(N__11365),
            .I(N__11362));
    InMux I__1780 (
            .O(N__11362),
            .I(N__11359));
    LocalMux I__1779 (
            .O(N__11359),
            .I(N__11355));
    CascadeMux I__1778 (
            .O(N__11358),
            .I(N__11349));
    Span4Mux_v I__1777 (
            .O(N__11355),
            .I(N__11340));
    InMux I__1776 (
            .O(N__11354),
            .I(N__11335));
    InMux I__1775 (
            .O(N__11353),
            .I(N__11335));
    InMux I__1774 (
            .O(N__11352),
            .I(N__11332));
    InMux I__1773 (
            .O(N__11349),
            .I(N__11325));
    InMux I__1772 (
            .O(N__11348),
            .I(N__11325));
    InMux I__1771 (
            .O(N__11347),
            .I(N__11325));
    InMux I__1770 (
            .O(N__11346),
            .I(N__11316));
    InMux I__1769 (
            .O(N__11345),
            .I(N__11316));
    InMux I__1768 (
            .O(N__11344),
            .I(N__11316));
    InMux I__1767 (
            .O(N__11343),
            .I(N__11316));
    Odrv4 I__1766 (
            .O(N__11340),
            .I(G_181));
    LocalMux I__1765 (
            .O(N__11335),
            .I(G_181));
    LocalMux I__1764 (
            .O(N__11332),
            .I(G_181));
    LocalMux I__1763 (
            .O(N__11325),
            .I(G_181));
    LocalMux I__1762 (
            .O(N__11316),
            .I(G_181));
    InMux I__1761 (
            .O(N__11305),
            .I(N__11302));
    LocalMux I__1760 (
            .O(N__11302),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ));
    CascadeMux I__1759 (
            .O(N__11299),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_ ));
    InMux I__1758 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__1757 (
            .O(N__11293),
            .I(N__11290));
    Odrv4 I__1756 (
            .O(N__11290),
            .I(\Lab_UT.didp.countrce1.q_5_3 ));
    CascadeMux I__1755 (
            .O(N__11287),
            .I(N__11284));
    InMux I__1754 (
            .O(N__11284),
            .I(N__11281));
    LocalMux I__1753 (
            .O(N__11281),
            .I(N__11278));
    Span4Mux_v I__1752 (
            .O(N__11278),
            .I(N__11275));
    Odrv4 I__1751 (
            .O(N__11275),
            .I(\Lab_UT.dispString.N_137 ));
    InMux I__1750 (
            .O(N__11272),
            .I(N__11269));
    LocalMux I__1749 (
            .O(N__11269),
            .I(N__11265));
    InMux I__1748 (
            .O(N__11268),
            .I(N__11262));
    Odrv4 I__1747 (
            .O(N__11265),
            .I(uu0_sec_clkD));
    LocalMux I__1746 (
            .O(N__11262),
            .I(uu0_sec_clkD));
    CascadeMux I__1745 (
            .O(N__11257),
            .I(\Lab_UT.dispString.N_143_cascade_ ));
    CascadeMux I__1744 (
            .O(N__11254),
            .I(N__11251));
    InMux I__1743 (
            .O(N__11251),
            .I(N__11247));
    InMux I__1742 (
            .O(N__11250),
            .I(N__11244));
    LocalMux I__1741 (
            .O(N__11247),
            .I(N__11239));
    LocalMux I__1740 (
            .O(N__11244),
            .I(N__11239));
    Span4Mux_h I__1739 (
            .O(N__11239),
            .I(N__11236));
    Odrv4 I__1738 (
            .O(N__11236),
            .I(\Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ));
    InMux I__1737 (
            .O(N__11233),
            .I(N__11230));
    LocalMux I__1736 (
            .O(N__11230),
            .I(N__11226));
    InMux I__1735 (
            .O(N__11229),
            .I(N__11223));
    Span4Mux_h I__1734 (
            .O(N__11226),
            .I(N__11220));
    LocalMux I__1733 (
            .O(N__11223),
            .I(N__11217));
    Odrv4 I__1732 (
            .O(N__11220),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    Odrv12 I__1731 (
            .O(N__11217),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__1730 (
            .O(N__11212),
            .I(N__11209));
    LocalMux I__1729 (
            .O(N__11209),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    InMux I__1728 (
            .O(N__11206),
            .I(N__11200));
    InMux I__1727 (
            .O(N__11205),
            .I(N__11200));
    LocalMux I__1726 (
            .O(N__11200),
            .I(N__11197));
    Sp12to4 I__1725 (
            .O(N__11197),
            .I(N__11194));
    Span12Mux_s3_v I__1724 (
            .O(N__11194),
            .I(N__11189));
    InMux I__1723 (
            .O(N__11193),
            .I(N__11184));
    InMux I__1722 (
            .O(N__11192),
            .I(N__11184));
    Odrv12 I__1721 (
            .O(N__11189),
            .I(\Lab_UT.didp.ce_12_1 ));
    LocalMux I__1720 (
            .O(N__11184),
            .I(\Lab_UT.didp.ce_12_1 ));
    CascadeMux I__1719 (
            .O(N__11179),
            .I(\Lab_UT.didp.ce_12_1_cascade_ ));
    CascadeMux I__1718 (
            .O(N__11176),
            .I(\Lab_UT.didp.ce_12_3_cascade_ ));
    CascadeMux I__1717 (
            .O(N__11173),
            .I(N__11170));
    InMux I__1716 (
            .O(N__11170),
            .I(N__11161));
    InMux I__1715 (
            .O(N__11169),
            .I(N__11161));
    InMux I__1714 (
            .O(N__11168),
            .I(N__11161));
    LocalMux I__1713 (
            .O(N__11161),
            .I(\Lab_UT.didp.countrce1.ce_12_1_1 ));
    CascadeMux I__1712 (
            .O(N__11158),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    CascadeMux I__1711 (
            .O(N__11155),
            .I(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ));
    CascadeMux I__1710 (
            .O(N__11152),
            .I(\Lab_UT.didp.countrce3.q_5_2_cascade_ ));
    InMux I__1709 (
            .O(N__11149),
            .I(N__11145));
    InMux I__1708 (
            .O(N__11148),
            .I(N__11142));
    LocalMux I__1707 (
            .O(N__11145),
            .I(N__11139));
    LocalMux I__1706 (
            .O(N__11142),
            .I(N__11136));
    Span4Mux_v I__1705 (
            .O(N__11139),
            .I(N__11132));
    Span4Mux_s2_v I__1704 (
            .O(N__11136),
            .I(N__11125));
    CascadeMux I__1703 (
            .O(N__11135),
            .I(N__11121));
    Span4Mux_h I__1702 (
            .O(N__11132),
            .I(N__11116));
    InMux I__1701 (
            .O(N__11131),
            .I(N__11113));
    CascadeMux I__1700 (
            .O(N__11130),
            .I(N__11107));
    CascadeMux I__1699 (
            .O(N__11129),
            .I(N__11104));
    CascadeMux I__1698 (
            .O(N__11128),
            .I(N__11101));
    Sp12to4 I__1697 (
            .O(N__11125),
            .I(N__11098));
    InMux I__1696 (
            .O(N__11124),
            .I(N__11089));
    InMux I__1695 (
            .O(N__11121),
            .I(N__11089));
    InMux I__1694 (
            .O(N__11120),
            .I(N__11089));
    InMux I__1693 (
            .O(N__11119),
            .I(N__11089));
    Span4Mux_v I__1692 (
            .O(N__11116),
            .I(N__11084));
    LocalMux I__1691 (
            .O(N__11113),
            .I(N__11084));
    InMux I__1690 (
            .O(N__11112),
            .I(N__11073));
    InMux I__1689 (
            .O(N__11111),
            .I(N__11073));
    InMux I__1688 (
            .O(N__11110),
            .I(N__11073));
    InMux I__1687 (
            .O(N__11107),
            .I(N__11073));
    InMux I__1686 (
            .O(N__11104),
            .I(N__11073));
    InMux I__1685 (
            .O(N__11101),
            .I(N__11070));
    Odrv12 I__1684 (
            .O(N__11098),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__1683 (
            .O(N__11089),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__1682 (
            .O(N__11084),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__1681 (
            .O(N__11073),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__1680 (
            .O(N__11070),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__1679 (
            .O(N__11059),
            .I(N__11056));
    LocalMux I__1678 (
            .O(N__11056),
            .I(\uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ));
    CascadeMux I__1677 (
            .O(N__11053),
            .I(N__11050));
    InMux I__1676 (
            .O(N__11050),
            .I(N__11044));
    InMux I__1675 (
            .O(N__11049),
            .I(N__11044));
    LocalMux I__1674 (
            .O(N__11044),
            .I(N__11041));
    Odrv4 I__1673 (
            .O(N__11041),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    CascadeMux I__1672 (
            .O(N__11038),
            .I(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ));
    InMux I__1671 (
            .O(N__11035),
            .I(N__11032));
    LocalMux I__1670 (
            .O(N__11032),
            .I(\uu2.bitmap_pmux_sn_i5_mux ));
    InMux I__1669 (
            .O(N__11029),
            .I(N__11025));
    InMux I__1668 (
            .O(N__11028),
            .I(N__11022));
    LocalMux I__1667 (
            .O(N__11025),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    LocalMux I__1666 (
            .O(N__11022),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    CascadeMux I__1665 (
            .O(N__11017),
            .I(\uu2.bitmap_pmux_sn_N_15_cascade_ ));
    InMux I__1664 (
            .O(N__11014),
            .I(N__11011));
    LocalMux I__1663 (
            .O(N__11011),
            .I(\uu2.N_401 ));
    InMux I__1662 (
            .O(N__11008),
            .I(N__11005));
    LocalMux I__1661 (
            .O(N__11005),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__1660 (
            .O(N__11002),
            .I(N__10984));
    InMux I__1659 (
            .O(N__11001),
            .I(N__10984));
    InMux I__1658 (
            .O(N__11000),
            .I(N__10984));
    InMux I__1657 (
            .O(N__10999),
            .I(N__10984));
    InMux I__1656 (
            .O(N__10998),
            .I(N__10984));
    InMux I__1655 (
            .O(N__10997),
            .I(N__10984));
    LocalMux I__1654 (
            .O(N__10984),
            .I(\uu2.un28_w_addr_user_i ));
    CascadeMux I__1653 (
            .O(N__10981),
            .I(N__10978));
    InMux I__1652 (
            .O(N__10978),
            .I(N__10974));
    InMux I__1651 (
            .O(N__10977),
            .I(N__10971));
    LocalMux I__1650 (
            .O(N__10974),
            .I(G_182));
    LocalMux I__1649 (
            .O(N__10971),
            .I(G_182));
    InMux I__1648 (
            .O(N__10966),
            .I(N__10957));
    InMux I__1647 (
            .O(N__10965),
            .I(N__10957));
    InMux I__1646 (
            .O(N__10964),
            .I(N__10957));
    LocalMux I__1645 (
            .O(N__10957),
            .I(G_183));
    CascadeMux I__1644 (
            .O(N__10954),
            .I(G_182_cascade_));
    InMux I__1643 (
            .O(N__10951),
            .I(N__10948));
    LocalMux I__1642 (
            .O(N__10948),
            .I(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ));
    CascadeMux I__1641 (
            .O(N__10945),
            .I(\Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ));
    InMux I__1640 (
            .O(N__10942),
            .I(N__10937));
    InMux I__1639 (
            .O(N__10941),
            .I(N__10932));
    InMux I__1638 (
            .O(N__10940),
            .I(N__10932));
    LocalMux I__1637 (
            .O(N__10937),
            .I(\Lab_UT.dictrl.alarmstateZ0Z8 ));
    LocalMux I__1636 (
            .O(N__10932),
            .I(\Lab_UT.dictrl.alarmstateZ0Z8 ));
    CascadeMux I__1635 (
            .O(N__10927),
            .I(\Lab_UT.dictrl.g1_0_4_0_cascade_ ));
    InMux I__1634 (
            .O(N__10924),
            .I(N__10921));
    LocalMux I__1633 (
            .O(N__10921),
            .I(\Lab_UT.dictrl.g1_0Z0Z_1 ));
    CascadeMux I__1632 (
            .O(N__10918),
            .I(\Lab_UT.dictrl.g0_5_4_0_cascade_ ));
    InMux I__1631 (
            .O(N__10915),
            .I(N__10911));
    InMux I__1630 (
            .O(N__10914),
            .I(N__10908));
    LocalMux I__1629 (
            .O(N__10911),
            .I(G_188));
    LocalMux I__1628 (
            .O(N__10908),
            .I(G_188));
    InMux I__1627 (
            .O(N__10903),
            .I(N__10900));
    LocalMux I__1626 (
            .O(N__10900),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_3 ));
    CascadeMux I__1625 (
            .O(N__10897),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_ ));
    InMux I__1624 (
            .O(N__10894),
            .I(N__10891));
    LocalMux I__1623 (
            .O(N__10891),
            .I(N__10888));
    Span4Mux_v I__1622 (
            .O(N__10888),
            .I(N__10883));
    InMux I__1621 (
            .O(N__10887),
            .I(N__10878));
    InMux I__1620 (
            .O(N__10886),
            .I(N__10878));
    Odrv4 I__1619 (
            .O(N__10883),
            .I(L3_tx_data_3));
    LocalMux I__1618 (
            .O(N__10878),
            .I(L3_tx_data_3));
    CascadeMux I__1617 (
            .O(N__10873),
            .I(G_186_cascade_));
    InMux I__1616 (
            .O(N__10870),
            .I(N__10864));
    InMux I__1615 (
            .O(N__10869),
            .I(N__10864));
    LocalMux I__1614 (
            .O(N__10864),
            .I(G_187));
    CascadeMux I__1613 (
            .O(N__10861),
            .I(G_187_cascade_));
    InMux I__1612 (
            .O(N__10858),
            .I(N__10855));
    LocalMux I__1611 (
            .O(N__10855),
            .I(\Lab_UT.dispString.dOutP_1_iv_i_1_4 ));
    CascadeMux I__1610 (
            .O(N__10852),
            .I(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ));
    IoInMux I__1609 (
            .O(N__10849),
            .I(N__10846));
    LocalMux I__1608 (
            .O(N__10846),
            .I(N__10842));
    SRMux I__1607 (
            .O(N__10845),
            .I(N__10839));
    IoSpan4Mux I__1606 (
            .O(N__10842),
            .I(N__10835));
    LocalMux I__1605 (
            .O(N__10839),
            .I(N__10832));
    CascadeMux I__1604 (
            .O(N__10838),
            .I(N__10829));
    Span4Mux_s1_v I__1603 (
            .O(N__10835),
            .I(N__10824));
    Span4Mux_h I__1602 (
            .O(N__10832),
            .I(N__10824));
    InMux I__1601 (
            .O(N__10829),
            .I(N__10821));
    Span4Mux_v I__1600 (
            .O(N__10824),
            .I(N__10816));
    LocalMux I__1599 (
            .O(N__10821),
            .I(N__10813));
    InMux I__1598 (
            .O(N__10820),
            .I(N__10810));
    InMux I__1597 (
            .O(N__10819),
            .I(N__10807));
    Odrv4 I__1596 (
            .O(N__10816),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1595 (
            .O(N__10813),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1594 (
            .O(N__10810),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1593 (
            .O(N__10807),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1592 (
            .O(N__10798),
            .I(\uu2.un1_w_user_lfZ0Z_4_cascade_ ));
    InMux I__1591 (
            .O(N__10795),
            .I(N__10789));
    InMux I__1590 (
            .O(N__10794),
            .I(N__10789));
    LocalMux I__1589 (
            .O(N__10789),
            .I(N__10786));
    Odrv12 I__1588 (
            .O(N__10786),
            .I(\uu2.un20_w_addr_userZ0Z_1 ));
    InMux I__1587 (
            .O(N__10783),
            .I(N__10780));
    LocalMux I__1586 (
            .O(N__10780),
            .I(N__10777));
    Span12Mux_s3_v I__1585 (
            .O(N__10777),
            .I(N__10772));
    InMux I__1584 (
            .O(N__10776),
            .I(N__10767));
    InMux I__1583 (
            .O(N__10775),
            .I(N__10767));
    Odrv12 I__1582 (
            .O(N__10772),
            .I(L3_tx_data_1));
    LocalMux I__1581 (
            .O(N__10767),
            .I(L3_tx_data_1));
    InMux I__1580 (
            .O(N__10762),
            .I(N__10759));
    LocalMux I__1579 (
            .O(N__10759),
            .I(N__10756));
    Span4Mux_s3_v I__1578 (
            .O(N__10756),
            .I(N__10751));
    InMux I__1577 (
            .O(N__10755),
            .I(N__10746));
    InMux I__1576 (
            .O(N__10754),
            .I(N__10746));
    Odrv4 I__1575 (
            .O(N__10751),
            .I(L3_tx_data_4));
    LocalMux I__1574 (
            .O(N__10746),
            .I(L3_tx_data_4));
    InMux I__1573 (
            .O(N__10741),
            .I(N__10737));
    CascadeMux I__1572 (
            .O(N__10740),
            .I(N__10734));
    LocalMux I__1571 (
            .O(N__10737),
            .I(N__10730));
    InMux I__1570 (
            .O(N__10734),
            .I(N__10727));
    InMux I__1569 (
            .O(N__10733),
            .I(N__10724));
    Odrv12 I__1568 (
            .O(N__10730),
            .I(L3_tx_data_6));
    LocalMux I__1567 (
            .O(N__10727),
            .I(L3_tx_data_6));
    LocalMux I__1566 (
            .O(N__10724),
            .I(L3_tx_data_6));
    InMux I__1565 (
            .O(N__10717),
            .I(N__10714));
    LocalMux I__1564 (
            .O(N__10714),
            .I(\uu2.un1_w_user_lfZ0Z_3 ));
    CascadeMux I__1563 (
            .O(N__10711),
            .I(N__10708));
    InMux I__1562 (
            .O(N__10708),
            .I(N__10705));
    LocalMux I__1561 (
            .O(N__10705),
            .I(N__10702));
    Odrv12 I__1560 (
            .O(N__10702),
            .I(\Lab_UT.dispString.N_140 ));
    InMux I__1559 (
            .O(N__10699),
            .I(N__10695));
    CascadeMux I__1558 (
            .O(N__10698),
            .I(N__10692));
    LocalMux I__1557 (
            .O(N__10695),
            .I(N__10689));
    InMux I__1556 (
            .O(N__10692),
            .I(N__10686));
    Span4Mux_v I__1555 (
            .O(N__10689),
            .I(N__10682));
    LocalMux I__1554 (
            .O(N__10686),
            .I(N__10679));
    InMux I__1553 (
            .O(N__10685),
            .I(N__10676));
    Odrv4 I__1552 (
            .O(N__10682),
            .I(L3_tx_data_5));
    Odrv4 I__1551 (
            .O(N__10679),
            .I(L3_tx_data_5));
    LocalMux I__1550 (
            .O(N__10676),
            .I(L3_tx_data_5));
    CascadeMux I__1549 (
            .O(N__10669),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ));
    InMux I__1548 (
            .O(N__10666),
            .I(N__10662));
    InMux I__1547 (
            .O(N__10665),
            .I(N__10659));
    LocalMux I__1546 (
            .O(N__10662),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    LocalMux I__1545 (
            .O(N__10659),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    InMux I__1544 (
            .O(N__10654),
            .I(N__10651));
    LocalMux I__1543 (
            .O(N__10651),
            .I(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ));
    InMux I__1542 (
            .O(N__10648),
            .I(N__10645));
    LocalMux I__1541 (
            .O(N__10645),
            .I(\uu2.w_addr_displaying_RNI0NG56Z0Z_4 ));
    InMux I__1540 (
            .O(N__10642),
            .I(N__10639));
    LocalMux I__1539 (
            .O(N__10639),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1538 (
            .O(N__10636),
            .I(N__10632));
    InMux I__1537 (
            .O(N__10635),
            .I(N__10629));
    LocalMux I__1536 (
            .O(N__10632),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    LocalMux I__1535 (
            .O(N__10629),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    InMux I__1534 (
            .O(N__10624),
            .I(N__10621));
    LocalMux I__1533 (
            .O(N__10621),
            .I(N__10618));
    Sp12to4 I__1532 (
            .O(N__10618),
            .I(N__10615));
    Span12Mux_s10_v I__1531 (
            .O(N__10615),
            .I(N__10612));
    Odrv12 I__1530 (
            .O(N__10612),
            .I(uart_RXD));
    SRMux I__1529 (
            .O(N__10609),
            .I(N__10605));
    CEMux I__1528 (
            .O(N__10608),
            .I(N__10602));
    LocalMux I__1527 (
            .O(N__10605),
            .I(N__10599));
    LocalMux I__1526 (
            .O(N__10602),
            .I(N__10596));
    Span4Mux_s3_h I__1525 (
            .O(N__10599),
            .I(N__10591));
    Span4Mux_s0_v I__1524 (
            .O(N__10596),
            .I(N__10591));
    Span4Mux_v I__1523 (
            .O(N__10591),
            .I(N__10588));
    Odrv4 I__1522 (
            .O(N__10588),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    InMux I__1521 (
            .O(N__10585),
            .I(N__10582));
    LocalMux I__1520 (
            .O(N__10582),
            .I(\uu2.w_addr_displaying_RNI03P31Z0Z_4 ));
    CascadeMux I__1519 (
            .O(N__10579),
            .I(\uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ));
    InMux I__1518 (
            .O(N__10576),
            .I(N__10573));
    LocalMux I__1517 (
            .O(N__10573),
            .I(\uu2.bitmap_pmux_sn_i7_mux_0 ));
    CascadeMux I__1516 (
            .O(N__10570),
            .I(\uu2.N_406_cascade_ ));
    InMux I__1515 (
            .O(N__10567),
            .I(N__10561));
    InMux I__1514 (
            .O(N__10566),
            .I(N__10561));
    LocalMux I__1513 (
            .O(N__10561),
            .I(\uu2.bitmap_pmux ));
    CascadeMux I__1512 (
            .O(N__10558),
            .I(\uu2.N_383_cascade_ ));
    CascadeMux I__1511 (
            .O(N__10555),
            .I(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ));
    InMux I__1510 (
            .O(N__10552),
            .I(N__10549));
    LocalMux I__1509 (
            .O(N__10549),
            .I(\uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ));
    InMux I__1508 (
            .O(N__10546),
            .I(N__10543));
    LocalMux I__1507 (
            .O(N__10543),
            .I(\uu2.bitmap_pmux_u_1 ));
    CascadeMux I__1506 (
            .O(N__10540),
            .I(\uu2.un28_w_addr_user_i_cascade_ ));
    CascadeMux I__1505 (
            .O(N__10537),
            .I(N__10533));
    CascadeMux I__1504 (
            .O(N__10536),
            .I(N__10530));
    InMux I__1503 (
            .O(N__10533),
            .I(N__10524));
    InMux I__1502 (
            .O(N__10530),
            .I(N__10524));
    InMux I__1501 (
            .O(N__10529),
            .I(N__10521));
    LocalMux I__1500 (
            .O(N__10524),
            .I(\uu2.un51_w_data_displaying_i_a2_1 ));
    LocalMux I__1499 (
            .O(N__10521),
            .I(\uu2.un51_w_data_displaying_i_a2_1 ));
    CascadeMux I__1498 (
            .O(N__10516),
            .I(\uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ));
    InMux I__1497 (
            .O(N__10513),
            .I(N__10507));
    InMux I__1496 (
            .O(N__10512),
            .I(N__10507));
    LocalMux I__1495 (
            .O(N__10507),
            .I(\uu2.w_data_displaying_2_i_a2_i_a3_2_0 ));
    CascadeMux I__1494 (
            .O(N__10504),
            .I(G_179_cascade_));
    InMux I__1493 (
            .O(N__10501),
            .I(N__10495));
    InMux I__1492 (
            .O(N__10500),
            .I(N__10488));
    InMux I__1491 (
            .O(N__10499),
            .I(N__10488));
    InMux I__1490 (
            .O(N__10498),
            .I(N__10488));
    LocalMux I__1489 (
            .O(N__10495),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    LocalMux I__1488 (
            .O(N__10488),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    CascadeMux I__1487 (
            .O(N__10483),
            .I(\Lab_UT.un1_idle_5_0_iclkZ0_cascade_ ));
    InMux I__1486 (
            .O(N__10480),
            .I(N__10476));
    InMux I__1485 (
            .O(N__10479),
            .I(N__10473));
    LocalMux I__1484 (
            .O(N__10476),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0 ));
    LocalMux I__1483 (
            .O(N__10473),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0 ));
    InMux I__1482 (
            .O(N__10468),
            .I(N__10464));
    InMux I__1481 (
            .O(N__10467),
            .I(N__10461));
    LocalMux I__1480 (
            .O(N__10464),
            .I(G_185));
    LocalMux I__1479 (
            .O(N__10461),
            .I(G_185));
    InMux I__1478 (
            .O(N__10456),
            .I(N__10453));
    LocalMux I__1477 (
            .O(N__10453),
            .I(N__10450));
    Span4Mux_h I__1476 (
            .O(N__10450),
            .I(N__10447));
    Odrv4 I__1475 (
            .O(N__10447),
            .I(vbuf_tx_data_6));
    InMux I__1474 (
            .O(N__10444),
            .I(N__10441));
    LocalMux I__1473 (
            .O(N__10441),
            .I(N__10438));
    Span4Mux_v I__1472 (
            .O(N__10438),
            .I(N__10435));
    Odrv4 I__1471 (
            .O(N__10435),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__1470 (
            .O(N__10432),
            .I(N__10429));
    LocalMux I__1469 (
            .O(N__10429),
            .I(N__10426));
    Odrv12 I__1468 (
            .O(N__10426),
            .I(vbuf_tx_data_7));
    InMux I__1467 (
            .O(N__10423),
            .I(N__10420));
    LocalMux I__1466 (
            .O(N__10420),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__1465 (
            .O(N__10417),
            .I(N__10414));
    InMux I__1464 (
            .O(N__10414),
            .I(N__10411));
    LocalMux I__1463 (
            .O(N__10411),
            .I(N__10408));
    Odrv4 I__1462 (
            .O(N__10408),
            .I(\uu2.mem0.w_addr_8 ));
    CEMux I__1461 (
            .O(N__10405),
            .I(N__10402));
    LocalMux I__1460 (
            .O(N__10402),
            .I(N__10399));
    Odrv4 I__1459 (
            .O(N__10399),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    CascadeMux I__1458 (
            .O(N__10396),
            .I(\Lab_UT.un1_idle_1_0_iclkZ0_cascade_ ));
    CascadeMux I__1457 (
            .O(N__10393),
            .I(\Lab_UT.dispString.N_117_cascade_ ));
    CascadeMux I__1456 (
            .O(N__10390),
            .I(G_180_cascade_));
    CascadeMux I__1455 (
            .O(N__10387),
            .I(G_181_cascade_));
    InMux I__1454 (
            .O(N__10384),
            .I(N__10381));
    LocalMux I__1453 (
            .O(N__10381),
            .I(G_180));
    CascadeMux I__1452 (
            .O(N__10378),
            .I(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ));
    InMux I__1451 (
            .O(N__10375),
            .I(N__10369));
    CascadeMux I__1450 (
            .O(N__10374),
            .I(N__10366));
    CascadeMux I__1449 (
            .O(N__10373),
            .I(N__10362));
    InMux I__1448 (
            .O(N__10372),
            .I(N__10359));
    LocalMux I__1447 (
            .O(N__10369),
            .I(N__10356));
    InMux I__1446 (
            .O(N__10366),
            .I(N__10351));
    InMux I__1445 (
            .O(N__10365),
            .I(N__10351));
    InMux I__1444 (
            .O(N__10362),
            .I(N__10348));
    LocalMux I__1443 (
            .O(N__10359),
            .I(\uu2.l_countZ0Z_1 ));
    Odrv4 I__1442 (
            .O(N__10356),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1441 (
            .O(N__10351),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1440 (
            .O(N__10348),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__1439 (
            .O(N__10339),
            .I(N__10334));
    InMux I__1438 (
            .O(N__10338),
            .I(N__10326));
    InMux I__1437 (
            .O(N__10337),
            .I(N__10326));
    LocalMux I__1436 (
            .O(N__10334),
            .I(N__10323));
    InMux I__1435 (
            .O(N__10333),
            .I(N__10320));
    InMux I__1434 (
            .O(N__10332),
            .I(N__10315));
    InMux I__1433 (
            .O(N__10331),
            .I(N__10315));
    LocalMux I__1432 (
            .O(N__10326),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__1431 (
            .O(N__10323),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1430 (
            .O(N__10320),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1429 (
            .O(N__10315),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__1428 (
            .O(N__10306),
            .I(N__10300));
    InMux I__1427 (
            .O(N__10305),
            .I(N__10300));
    LocalMux I__1426 (
            .O(N__10300),
            .I(N__10297));
    Odrv12 I__1425 (
            .O(N__10297),
            .I(\uu2.un284_ci ));
    CascadeMux I__1424 (
            .O(N__10294),
            .I(\Lab_UT.didp.countrce1.q_5_0_cascade_ ));
    CEMux I__1423 (
            .O(N__10291),
            .I(N__10287));
    CEMux I__1422 (
            .O(N__10290),
            .I(N__10284));
    LocalMux I__1421 (
            .O(N__10287),
            .I(N__10281));
    LocalMux I__1420 (
            .O(N__10284),
            .I(N__10278));
    Span4Mux_v I__1419 (
            .O(N__10281),
            .I(N__10275));
    Odrv12 I__1418 (
            .O(N__10278),
            .I(\Lab_UT.didp.regrce3.LdAMones_0 ));
    Odrv4 I__1417 (
            .O(N__10275),
            .I(\Lab_UT.didp.regrce3.LdAMones_0 ));
    InMux I__1416 (
            .O(N__10270),
            .I(N__10267));
    LocalMux I__1415 (
            .O(N__10267),
            .I(G_184));
    CascadeMux I__1414 (
            .O(N__10264),
            .I(G_184_cascade_));
    CascadeMux I__1413 (
            .O(N__10261),
            .I(N__10256));
    InMux I__1412 (
            .O(N__10260),
            .I(N__10248));
    InMux I__1411 (
            .O(N__10259),
            .I(N__10248));
    InMux I__1410 (
            .O(N__10256),
            .I(N__10245));
    InMux I__1409 (
            .O(N__10255),
            .I(N__10238));
    InMux I__1408 (
            .O(N__10254),
            .I(N__10238));
    InMux I__1407 (
            .O(N__10253),
            .I(N__10238));
    LocalMux I__1406 (
            .O(N__10248),
            .I(N__10235));
    LocalMux I__1405 (
            .O(N__10245),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1404 (
            .O(N__10238),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__1403 (
            .O(N__10235),
            .I(\uu2.r_addrZ0Z_0 ));
    CEMux I__1402 (
            .O(N__10228),
            .I(N__10225));
    LocalMux I__1401 (
            .O(N__10225),
            .I(N__10222));
    Odrv12 I__1400 (
            .O(N__10222),
            .I(\uu2.trig_rd_is_det_0 ));
    InMux I__1399 (
            .O(N__10219),
            .I(N__10216));
    LocalMux I__1398 (
            .O(N__10216),
            .I(N__10213));
    Span4Mux_s0_v I__1397 (
            .O(N__10213),
            .I(N__10210));
    Odrv4 I__1396 (
            .O(N__10210),
            .I(\uu2.mem0.w_data_2 ));
    CascadeMux I__1395 (
            .O(N__10207),
            .I(N__10201));
    InMux I__1394 (
            .O(N__10206),
            .I(N__10198));
    InMux I__1393 (
            .O(N__10205),
            .I(N__10192));
    InMux I__1392 (
            .O(N__10204),
            .I(N__10192));
    InMux I__1391 (
            .O(N__10201),
            .I(N__10189));
    LocalMux I__1390 (
            .O(N__10198),
            .I(N__10186));
    InMux I__1389 (
            .O(N__10197),
            .I(N__10183));
    LocalMux I__1388 (
            .O(N__10192),
            .I(N__10180));
    LocalMux I__1387 (
            .O(N__10189),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1386 (
            .O(N__10186),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1385 (
            .O(N__10183),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1384 (
            .O(N__10180),
            .I(\uu2.r_addrZ0Z_4 ));
    CascadeMux I__1383 (
            .O(N__10171),
            .I(N__10168));
    InMux I__1382 (
            .O(N__10168),
            .I(N__10162));
    InMux I__1381 (
            .O(N__10167),
            .I(N__10159));
    InMux I__1380 (
            .O(N__10166),
            .I(N__10156));
    InMux I__1379 (
            .O(N__10165),
            .I(N__10153));
    LocalMux I__1378 (
            .O(N__10162),
            .I(N__10146));
    LocalMux I__1377 (
            .O(N__10159),
            .I(N__10146));
    LocalMux I__1376 (
            .O(N__10156),
            .I(N__10146));
    LocalMux I__1375 (
            .O(N__10153),
            .I(\uu2.un404_ci_0 ));
    Odrv12 I__1374 (
            .O(N__10146),
            .I(\uu2.un404_ci_0 ));
    InMux I__1373 (
            .O(N__10141),
            .I(N__10133));
    InMux I__1372 (
            .O(N__10140),
            .I(N__10122));
    InMux I__1371 (
            .O(N__10139),
            .I(N__10122));
    InMux I__1370 (
            .O(N__10138),
            .I(N__10122));
    InMux I__1369 (
            .O(N__10137),
            .I(N__10122));
    InMux I__1368 (
            .O(N__10136),
            .I(N__10122));
    LocalMux I__1367 (
            .O(N__10133),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__1366 (
            .O(N__10122),
            .I(\uu2.trig_rd_is_det ));
    InMux I__1365 (
            .O(N__10117),
            .I(N__10113));
    CascadeMux I__1364 (
            .O(N__10116),
            .I(N__10110));
    LocalMux I__1363 (
            .O(N__10113),
            .I(N__10107));
    InMux I__1362 (
            .O(N__10110),
            .I(N__10104));
    Span4Mux_s0_v I__1361 (
            .O(N__10107),
            .I(N__10097));
    LocalMux I__1360 (
            .O(N__10104),
            .I(N__10097));
    InMux I__1359 (
            .O(N__10103),
            .I(N__10094));
    CascadeMux I__1358 (
            .O(N__10102),
            .I(N__10091));
    Span4Mux_v I__1357 (
            .O(N__10097),
            .I(N__10086));
    LocalMux I__1356 (
            .O(N__10094),
            .I(N__10086));
    InMux I__1355 (
            .O(N__10091),
            .I(N__10083));
    Span4Mux_s0_v I__1354 (
            .O(N__10086),
            .I(N__10080));
    LocalMux I__1353 (
            .O(N__10083),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__1352 (
            .O(N__10080),
            .I(\uu2.r_addrZ0Z_5 ));
    InMux I__1351 (
            .O(N__10075),
            .I(N__10072));
    LocalMux I__1350 (
            .O(N__10072),
            .I(N__10065));
    InMux I__1349 (
            .O(N__10071),
            .I(N__10056));
    InMux I__1348 (
            .O(N__10070),
            .I(N__10056));
    InMux I__1347 (
            .O(N__10069),
            .I(N__10056));
    InMux I__1346 (
            .O(N__10068),
            .I(N__10056));
    Odrv4 I__1345 (
            .O(N__10065),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__1344 (
            .O(N__10056),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__1343 (
            .O(N__10051),
            .I(N__10048));
    InMux I__1342 (
            .O(N__10048),
            .I(N__10045));
    LocalMux I__1341 (
            .O(N__10045),
            .I(N__10041));
    InMux I__1340 (
            .O(N__10044),
            .I(N__10038));
    Odrv12 I__1339 (
            .O(N__10041),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    LocalMux I__1338 (
            .O(N__10038),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    InMux I__1337 (
            .O(N__10033),
            .I(N__10030));
    LocalMux I__1336 (
            .O(N__10030),
            .I(N__10027));
    Span4Mux_h I__1335 (
            .O(N__10027),
            .I(N__10020));
    InMux I__1334 (
            .O(N__10026),
            .I(N__10011));
    InMux I__1333 (
            .O(N__10025),
            .I(N__10011));
    InMux I__1332 (
            .O(N__10024),
            .I(N__10011));
    InMux I__1331 (
            .O(N__10023),
            .I(N__10011));
    Odrv4 I__1330 (
            .O(N__10020),
            .I(\uu2.un306_ci ));
    LocalMux I__1329 (
            .O(N__10011),
            .I(\uu2.un306_ci ));
    InMux I__1328 (
            .O(N__10006),
            .I(N__10002));
    InMux I__1327 (
            .O(N__10005),
            .I(N__9998));
    LocalMux I__1326 (
            .O(N__10002),
            .I(N__9995));
    InMux I__1325 (
            .O(N__10001),
            .I(N__9992));
    LocalMux I__1324 (
            .O(N__9998),
            .I(N__9989));
    Span4Mux_s3_h I__1323 (
            .O(N__9995),
            .I(N__9986));
    LocalMux I__1322 (
            .O(N__9992),
            .I(\uu2.l_countZ0Z_7 ));
    Odrv12 I__1321 (
            .O(N__9989),
            .I(\uu2.l_countZ0Z_7 ));
    Odrv4 I__1320 (
            .O(N__9986),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__1319 (
            .O(N__9979),
            .I(N__9976));
    LocalMux I__1318 (
            .O(N__9976),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1317 (
            .O(N__9973),
            .I(N__9970));
    LocalMux I__1316 (
            .O(N__9970),
            .I(\uu2.N_34 ));
    CascadeMux I__1315 (
            .O(N__9967),
            .I(\uu2.N_34_cascade_ ));
    InMux I__1314 (
            .O(N__9964),
            .I(N__9961));
    LocalMux I__1313 (
            .O(N__9961),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1312 (
            .O(N__9958),
            .I(N__9955));
    LocalMux I__1311 (
            .O(N__9955),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__1310 (
            .O(N__9952),
            .I(N__9949));
    LocalMux I__1309 (
            .O(N__9949),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1308 (
            .O(N__9946),
            .I(N__9940));
    InMux I__1307 (
            .O(N__9945),
            .I(N__9940));
    LocalMux I__1306 (
            .O(N__9940),
            .I(\uu2.N_31 ));
    CascadeMux I__1305 (
            .O(N__9937),
            .I(\uu2.N_31_cascade_ ));
    InMux I__1304 (
            .O(N__9934),
            .I(N__9931));
    LocalMux I__1303 (
            .O(N__9931),
            .I(\uu2.mem0.w_data_0 ));
    CascadeMux I__1302 (
            .O(N__9928),
            .I(N__9923));
    InMux I__1301 (
            .O(N__9927),
            .I(N__9917));
    InMux I__1300 (
            .O(N__9926),
            .I(N__9917));
    InMux I__1299 (
            .O(N__9923),
            .I(N__9914));
    InMux I__1298 (
            .O(N__9922),
            .I(N__9911));
    LocalMux I__1297 (
            .O(N__9917),
            .I(N__9908));
    LocalMux I__1296 (
            .O(N__9914),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1295 (
            .O(N__9911),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__1294 (
            .O(N__9908),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1293 (
            .O(N__9901),
            .I(N__9897));
    CascadeMux I__1292 (
            .O(N__9900),
            .I(N__9892));
    InMux I__1291 (
            .O(N__9897),
            .I(N__9888));
    InMux I__1290 (
            .O(N__9896),
            .I(N__9883));
    InMux I__1289 (
            .O(N__9895),
            .I(N__9883));
    InMux I__1288 (
            .O(N__9892),
            .I(N__9878));
    InMux I__1287 (
            .O(N__9891),
            .I(N__9878));
    LocalMux I__1286 (
            .O(N__9888),
            .I(N__9873));
    LocalMux I__1285 (
            .O(N__9883),
            .I(N__9873));
    LocalMux I__1284 (
            .O(N__9878),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv4 I__1283 (
            .O(N__9873),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1282 (
            .O(N__9868),
            .I(\uu2.vbuf_raddr.un448_ci_0_cascade_ ));
    CascadeMux I__1281 (
            .O(N__9865),
            .I(N__9862));
    InMux I__1280 (
            .O(N__9862),
            .I(N__9858));
    InMux I__1279 (
            .O(N__9861),
            .I(N__9855));
    LocalMux I__1278 (
            .O(N__9858),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1277 (
            .O(N__9855),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__1276 (
            .O(N__9850),
            .I(N__9847));
    InMux I__1275 (
            .O(N__9847),
            .I(N__9842));
    InMux I__1274 (
            .O(N__9846),
            .I(N__9837));
    InMux I__1273 (
            .O(N__9845),
            .I(N__9837));
    LocalMux I__1272 (
            .O(N__9842),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1271 (
            .O(N__9837),
            .I(\uu2.r_addrZ0Z_7 ));
    CascadeMux I__1270 (
            .O(N__9832),
            .I(N__9827));
    CascadeMux I__1269 (
            .O(N__9831),
            .I(N__9824));
    CascadeMux I__1268 (
            .O(N__9830),
            .I(N__9821));
    InMux I__1267 (
            .O(N__9827),
            .I(N__9818));
    InMux I__1266 (
            .O(N__9824),
            .I(N__9813));
    InMux I__1265 (
            .O(N__9821),
            .I(N__9813));
    LocalMux I__1264 (
            .O(N__9818),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1263 (
            .O(N__9813),
            .I(\uu2.r_addrZ0Z_3 ));
    CascadeMux I__1262 (
            .O(N__9808),
            .I(\uu2.un404_ci_0_cascade_ ));
    CascadeMux I__1261 (
            .O(N__9805),
            .I(N__9802));
    InMux I__1260 (
            .O(N__9802),
            .I(N__9796));
    InMux I__1259 (
            .O(N__9801),
            .I(N__9789));
    InMux I__1258 (
            .O(N__9800),
            .I(N__9789));
    InMux I__1257 (
            .O(N__9799),
            .I(N__9789));
    LocalMux I__1256 (
            .O(N__9796),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1255 (
            .O(N__9789),
            .I(\uu2.r_addrZ0Z_6 ));
    InMux I__1254 (
            .O(N__9784),
            .I(N__9778));
    InMux I__1253 (
            .O(N__9783),
            .I(N__9778));
    LocalMux I__1252 (
            .O(N__9778),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    InMux I__1251 (
            .O(N__9775),
            .I(N__9772));
    LocalMux I__1250 (
            .O(N__9772),
            .I(\uu2.mem0.w_data_6 ));
    CEMux I__1249 (
            .O(N__9769),
            .I(N__9763));
    CEMux I__1248 (
            .O(N__9768),
            .I(N__9760));
    CEMux I__1247 (
            .O(N__9767),
            .I(N__9757));
    CEMux I__1246 (
            .O(N__9766),
            .I(N__9754));
    LocalMux I__1245 (
            .O(N__9763),
            .I(N__9749));
    LocalMux I__1244 (
            .O(N__9760),
            .I(N__9749));
    LocalMux I__1243 (
            .O(N__9757),
            .I(N__9746));
    LocalMux I__1242 (
            .O(N__9754),
            .I(N__9743));
    Odrv4 I__1241 (
            .O(N__9749),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv12 I__1240 (
            .O(N__9746),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__1239 (
            .O(N__9743),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__1238 (
            .O(N__9736),
            .I(N__9731));
    InMux I__1237 (
            .O(N__9735),
            .I(N__9726));
    InMux I__1236 (
            .O(N__9734),
            .I(N__9726));
    LocalMux I__1235 (
            .O(N__9731),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1234 (
            .O(N__9726),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__1233 (
            .O(N__9721),
            .I(N__9717));
    CascadeMux I__1232 (
            .O(N__9720),
            .I(N__9713));
    InMux I__1231 (
            .O(N__9717),
            .I(N__9709));
    InMux I__1230 (
            .O(N__9716),
            .I(N__9702));
    InMux I__1229 (
            .O(N__9713),
            .I(N__9702));
    InMux I__1228 (
            .O(N__9712),
            .I(N__9702));
    LocalMux I__1227 (
            .O(N__9709),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1226 (
            .O(N__9702),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__1225 (
            .O(N__9697),
            .I(N__9692));
    InMux I__1224 (
            .O(N__9696),
            .I(N__9687));
    InMux I__1223 (
            .O(N__9695),
            .I(N__9687));
    LocalMux I__1222 (
            .O(N__9692),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1221 (
            .O(N__9687),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1220 (
            .O(N__9682),
            .I(N__9679));
    LocalMux I__1219 (
            .O(N__9679),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__1218 (
            .O(N__9676),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1217 (
            .O(N__9673),
            .I(N__9669));
    InMux I__1216 (
            .O(N__9672),
            .I(N__9666));
    LocalMux I__1215 (
            .O(N__9669),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__1214 (
            .O(N__9666),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1213 (
            .O(N__9661),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1212 (
            .O(N__9658),
            .I(N__9653));
    InMux I__1211 (
            .O(N__9657),
            .I(N__9648));
    InMux I__1210 (
            .O(N__9656),
            .I(N__9648));
    LocalMux I__1209 (
            .O(N__9653),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1208 (
            .O(N__9648),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1207 (
            .O(N__9643),
            .I(N__9640));
    InMux I__1206 (
            .O(N__9640),
            .I(N__9637));
    LocalMux I__1205 (
            .O(N__9637),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__1204 (
            .O(N__9634),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    CascadeMux I__1203 (
            .O(N__9631),
            .I(N__9625));
    InMux I__1202 (
            .O(N__9630),
            .I(N__9622));
    InMux I__1201 (
            .O(N__9629),
            .I(N__9615));
    InMux I__1200 (
            .O(N__9628),
            .I(N__9615));
    InMux I__1199 (
            .O(N__9625),
            .I(N__9615));
    LocalMux I__1198 (
            .O(N__9622),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1197 (
            .O(N__9615),
            .I(\buart.Z_rx.ser_clk ));
    InMux I__1196 (
            .O(N__9610),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__1195 (
            .O(N__9607),
            .I(N__9603));
    CascadeMux I__1194 (
            .O(N__9606),
            .I(N__9600));
    InMux I__1193 (
            .O(N__9603),
            .I(N__9597));
    InMux I__1192 (
            .O(N__9600),
            .I(N__9594));
    LocalMux I__1191 (
            .O(N__9597),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__1190 (
            .O(N__9594),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__1189 (
            .O(N__9589),
            .I(N__9582));
    InMux I__1188 (
            .O(N__9588),
            .I(N__9582));
    InMux I__1187 (
            .O(N__9587),
            .I(N__9579));
    LocalMux I__1186 (
            .O(N__9582),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__1185 (
            .O(N__9579),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__1184 (
            .O(N__9574),
            .I(N__9571));
    InMux I__1183 (
            .O(N__9571),
            .I(N__9561));
    InMux I__1182 (
            .O(N__9570),
            .I(N__9561));
    InMux I__1181 (
            .O(N__9569),
            .I(N__9561));
    InMux I__1180 (
            .O(N__9568),
            .I(N__9558));
    LocalMux I__1179 (
            .O(N__9561),
            .I(\resetGen.reset_countZ0Z_0 ));
    LocalMux I__1178 (
            .O(N__9558),
            .I(\resetGen.reset_countZ0Z_0 ));
    CascadeMux I__1177 (
            .O(N__9553),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__1176 (
            .O(N__9550),
            .I(N__9546));
    InMux I__1175 (
            .O(N__9549),
            .I(N__9543));
    LocalMux I__1174 (
            .O(N__9546),
            .I(\resetGen.reset_countZ0Z_3 ));
    LocalMux I__1173 (
            .O(N__9543),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__1172 (
            .O(N__9538),
            .I(N__9531));
    InMux I__1171 (
            .O(N__9537),
            .I(N__9521));
    InMux I__1170 (
            .O(N__9536),
            .I(N__9521));
    InMux I__1169 (
            .O(N__9535),
            .I(N__9521));
    InMux I__1168 (
            .O(N__9534),
            .I(N__9521));
    InMux I__1167 (
            .O(N__9531),
            .I(N__9516));
    InMux I__1166 (
            .O(N__9530),
            .I(N__9516));
    LocalMux I__1165 (
            .O(N__9521),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__1164 (
            .O(N__9516),
            .I(\resetGen.reset_countZ0Z_4 ));
    InMux I__1163 (
            .O(N__9511),
            .I(N__9505));
    InMux I__1162 (
            .O(N__9510),
            .I(N__9505));
    LocalMux I__1161 (
            .O(N__9505),
            .I(N__9502));
    Odrv4 I__1160 (
            .O(N__9502),
            .I(\resetGen.un241_ci ));
    CascadeMux I__1159 (
            .O(N__9499),
            .I(N__9496));
    InMux I__1158 (
            .O(N__9496),
            .I(N__9489));
    InMux I__1157 (
            .O(N__9495),
            .I(N__9489));
    InMux I__1156 (
            .O(N__9494),
            .I(N__9486));
    LocalMux I__1155 (
            .O(N__9489),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1154 (
            .O(N__9486),
            .I(\resetGen.reset_countZ0Z_2 ));
    CascadeMux I__1153 (
            .O(N__9481),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    InMux I__1152 (
            .O(N__9478),
            .I(N__9475));
    LocalMux I__1151 (
            .O(N__9475),
            .I(N__9472));
    Odrv4 I__1150 (
            .O(N__9472),
            .I(\buart.Z_rx.un1_sample_0 ));
    CascadeMux I__1149 (
            .O(N__9469),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    CascadeMux I__1148 (
            .O(N__9466),
            .I(N__9462));
    InMux I__1147 (
            .O(N__9465),
            .I(N__9458));
    InMux I__1146 (
            .O(N__9462),
            .I(N__9455));
    InMux I__1145 (
            .O(N__9461),
            .I(N__9450));
    LocalMux I__1144 (
            .O(N__9458),
            .I(N__9445));
    LocalMux I__1143 (
            .O(N__9455),
            .I(N__9445));
    InMux I__1142 (
            .O(N__9454),
            .I(N__9440));
    InMux I__1141 (
            .O(N__9453),
            .I(N__9440));
    LocalMux I__1140 (
            .O(N__9450),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv4 I__1139 (
            .O(N__9445),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__1138 (
            .O(N__9440),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    IoInMux I__1137 (
            .O(N__9433),
            .I(N__9430));
    LocalMux I__1136 (
            .O(N__9430),
            .I(N__9427));
    Span12Mux_s4_v I__1135 (
            .O(N__9427),
            .I(N__9424));
    Odrv12 I__1134 (
            .O(N__9424),
            .I(\buart.Z_rx.sample ));
    CascadeMux I__1133 (
            .O(N__9421),
            .I(N__9418));
    InMux I__1132 (
            .O(N__9418),
            .I(N__9415));
    LocalMux I__1131 (
            .O(N__9415),
            .I(N__9412));
    Odrv4 I__1130 (
            .O(N__9412),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    CascadeMux I__1129 (
            .O(N__9409),
            .I(N__9406));
    InMux I__1128 (
            .O(N__9406),
            .I(N__9402));
    InMux I__1127 (
            .O(N__9405),
            .I(N__9396));
    LocalMux I__1126 (
            .O(N__9402),
            .I(N__9393));
    InMux I__1125 (
            .O(N__9401),
            .I(N__9386));
    InMux I__1124 (
            .O(N__9400),
            .I(N__9386));
    InMux I__1123 (
            .O(N__9399),
            .I(N__9386));
    LocalMux I__1122 (
            .O(N__9396),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    Odrv4 I__1121 (
            .O(N__9393),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1120 (
            .O(N__9386),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    InMux I__1119 (
            .O(N__9379),
            .I(N__9374));
    InMux I__1118 (
            .O(N__9378),
            .I(N__9368));
    InMux I__1117 (
            .O(N__9377),
            .I(N__9368));
    LocalMux I__1116 (
            .O(N__9374),
            .I(N__9365));
    InMux I__1115 (
            .O(N__9373),
            .I(N__9362));
    LocalMux I__1114 (
            .O(N__9368),
            .I(\buart.Z_rx.N_27_0_i ));
    Odrv4 I__1113 (
            .O(N__9365),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1112 (
            .O(N__9362),
            .I(\buart.Z_rx.N_27_0_i ));
    InMux I__1111 (
            .O(N__9355),
            .I(N__9352));
    LocalMux I__1110 (
            .O(N__9352),
            .I(\uu0.delay_lineZ0Z_1 ));
    InMux I__1109 (
            .O(N__9349),
            .I(N__9345));
    InMux I__1108 (
            .O(N__9348),
            .I(N__9342));
    LocalMux I__1107 (
            .O(N__9345),
            .I(\uu0.delay_lineZ0Z_0 ));
    LocalMux I__1106 (
            .O(N__9342),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__1105 (
            .O(N__9337),
            .I(N__9333));
    InMux I__1104 (
            .O(N__9336),
            .I(N__9327));
    LocalMux I__1103 (
            .O(N__9333),
            .I(N__9317));
    InMux I__1102 (
            .O(N__9332),
            .I(N__9310));
    InMux I__1101 (
            .O(N__9331),
            .I(N__9310));
    InMux I__1100 (
            .O(N__9330),
            .I(N__9310));
    LocalMux I__1099 (
            .O(N__9327),
            .I(N__9307));
    InMux I__1098 (
            .O(N__9326),
            .I(N__9299));
    InMux I__1097 (
            .O(N__9325),
            .I(N__9299));
    InMux I__1096 (
            .O(N__9324),
            .I(N__9299));
    InMux I__1095 (
            .O(N__9323),
            .I(N__9296));
    InMux I__1094 (
            .O(N__9322),
            .I(N__9293));
    InMux I__1093 (
            .O(N__9321),
            .I(N__9290));
    InMux I__1092 (
            .O(N__9320),
            .I(N__9287));
    Span4Mux_v I__1091 (
            .O(N__9317),
            .I(N__9284));
    LocalMux I__1090 (
            .O(N__9310),
            .I(N__9279));
    Span4Mux_v I__1089 (
            .O(N__9307),
            .I(N__9279));
    InMux I__1088 (
            .O(N__9306),
            .I(N__9276));
    LocalMux I__1087 (
            .O(N__9299),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1086 (
            .O(N__9296),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1085 (
            .O(N__9293),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1084 (
            .O(N__9290),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1083 (
            .O(N__9287),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1082 (
            .O(N__9284),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1081 (
            .O(N__9279),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1080 (
            .O(N__9276),
            .I(\uu0.un4_l_count_0 ));
    IoInMux I__1079 (
            .O(N__9259),
            .I(N__9256));
    LocalMux I__1078 (
            .O(N__9256),
            .I(N__9253));
    Span4Mux_s1_h I__1077 (
            .O(N__9253),
            .I(N__9250));
    Odrv4 I__1076 (
            .O(N__9250),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__1075 (
            .O(N__9247),
            .I(N__9244));
    InMux I__1074 (
            .O(N__9244),
            .I(N__9241));
    LocalMux I__1073 (
            .O(N__9241),
            .I(N__9238));
    Span12Mux_s9_v I__1072 (
            .O(N__9238),
            .I(N__9235));
    Odrv12 I__1071 (
            .O(N__9235),
            .I(\uu2.mem0.w_addr_0 ));
    InMux I__1070 (
            .O(N__9232),
            .I(N__9229));
    LocalMux I__1069 (
            .O(N__9229),
            .I(\resetGen.reset_count_2_0_4 ));
    CascadeMux I__1068 (
            .O(N__9226),
            .I(N__9223));
    InMux I__1067 (
            .O(N__9223),
            .I(N__9220));
    LocalMux I__1066 (
            .O(N__9220),
            .I(\uu0.un99_ci_0 ));
    InMux I__1065 (
            .O(N__9217),
            .I(N__9212));
    InMux I__1064 (
            .O(N__9216),
            .I(N__9207));
    InMux I__1063 (
            .O(N__9215),
            .I(N__9207));
    LocalMux I__1062 (
            .O(N__9212),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__1061 (
            .O(N__9207),
            .I(\uu0.l_countZ0Z_7 ));
    InMux I__1060 (
            .O(N__9202),
            .I(N__9199));
    LocalMux I__1059 (
            .O(N__9199),
            .I(\uu0.un44_ci ));
    CascadeMux I__1058 (
            .O(N__9196),
            .I(\uu0.un44_ci_cascade_ ));
    InMux I__1057 (
            .O(N__9193),
            .I(N__9188));
    InMux I__1056 (
            .O(N__9192),
            .I(N__9183));
    InMux I__1055 (
            .O(N__9191),
            .I(N__9183));
    LocalMux I__1054 (
            .O(N__9188),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__1053 (
            .O(N__9183),
            .I(\uu0.l_countZ0Z_3 ));
    CascadeMux I__1052 (
            .O(N__9178),
            .I(N__9175));
    InMux I__1051 (
            .O(N__9175),
            .I(N__9172));
    LocalMux I__1050 (
            .O(N__9172),
            .I(N__9166));
    InMux I__1049 (
            .O(N__9171),
            .I(N__9161));
    InMux I__1048 (
            .O(N__9170),
            .I(N__9161));
    InMux I__1047 (
            .O(N__9169),
            .I(N__9158));
    Odrv4 I__1046 (
            .O(N__9166),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__1045 (
            .O(N__9161),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__1044 (
            .O(N__9158),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__1043 (
            .O(N__9151),
            .I(N__9144));
    CascadeMux I__1042 (
            .O(N__9150),
            .I(N__9141));
    InMux I__1041 (
            .O(N__9149),
            .I(N__9132));
    InMux I__1040 (
            .O(N__9148),
            .I(N__9132));
    InMux I__1039 (
            .O(N__9147),
            .I(N__9132));
    InMux I__1038 (
            .O(N__9144),
            .I(N__9132));
    InMux I__1037 (
            .O(N__9141),
            .I(N__9129));
    LocalMux I__1036 (
            .O(N__9132),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__1035 (
            .O(N__9129),
            .I(\uu0.l_countZ0Z_0 ));
    InMux I__1034 (
            .O(N__9124),
            .I(N__9114));
    InMux I__1033 (
            .O(N__9123),
            .I(N__9114));
    InMux I__1032 (
            .O(N__9122),
            .I(N__9114));
    InMux I__1031 (
            .O(N__9121),
            .I(N__9111));
    LocalMux I__1030 (
            .O(N__9114),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__1029 (
            .O(N__9111),
            .I(\uu0.l_countZ0Z_1 ));
    CascadeMux I__1028 (
            .O(N__9106),
            .I(\uu0.un66_ci_cascade_ ));
    CascadeMux I__1027 (
            .O(N__9103),
            .I(N__9100));
    InMux I__1026 (
            .O(N__9100),
            .I(N__9092));
    InMux I__1025 (
            .O(N__9099),
            .I(N__9092));
    InMux I__1024 (
            .O(N__9098),
            .I(N__9089));
    InMux I__1023 (
            .O(N__9097),
            .I(N__9086));
    LocalMux I__1022 (
            .O(N__9092),
            .I(N__9083));
    LocalMux I__1021 (
            .O(N__9089),
            .I(\uu0.un66_ci ));
    LocalMux I__1020 (
            .O(N__9086),
            .I(\uu0.un66_ci ));
    Odrv4 I__1019 (
            .O(N__9083),
            .I(\uu0.un66_ci ));
    CEMux I__1018 (
            .O(N__9076),
            .I(N__9064));
    CEMux I__1017 (
            .O(N__9075),
            .I(N__9064));
    CEMux I__1016 (
            .O(N__9074),
            .I(N__9064));
    CEMux I__1015 (
            .O(N__9073),
            .I(N__9064));
    GlobalMux I__1014 (
            .O(N__9064),
            .I(N__9061));
    gio2CtrlBuf I__1013 (
            .O(N__9061),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__1012 (
            .O(N__9058),
            .I(N__9055));
    InMux I__1011 (
            .O(N__9055),
            .I(N__9045));
    InMux I__1010 (
            .O(N__9054),
            .I(N__9045));
    InMux I__1009 (
            .O(N__9053),
            .I(N__9045));
    InMux I__1008 (
            .O(N__9052),
            .I(N__9042));
    LocalMux I__1007 (
            .O(N__9045),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__1006 (
            .O(N__9042),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__1005 (
            .O(N__9037),
            .I(N__9030));
    InMux I__1004 (
            .O(N__9036),
            .I(N__9030));
    InMux I__1003 (
            .O(N__9035),
            .I(N__9027));
    LocalMux I__1002 (
            .O(N__9030),
            .I(\uu0.l_countZ0Z_5 ));
    LocalMux I__1001 (
            .O(N__9027),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__1000 (
            .O(N__9022),
            .I(N__9017));
    InMux I__999 (
            .O(N__9021),
            .I(N__9010));
    InMux I__998 (
            .O(N__9020),
            .I(N__9010));
    InMux I__997 (
            .O(N__9017),
            .I(N__9010));
    LocalMux I__996 (
            .O(N__9010),
            .I(N__9007));
    Odrv4 I__995 (
            .O(N__9007),
            .I(\uu0.un88_ci_3 ));
    InMux I__994 (
            .O(N__9004),
            .I(N__9001));
    LocalMux I__993 (
            .O(N__9001),
            .I(N__8998));
    Odrv4 I__992 (
            .O(N__8998),
            .I(\uu0.un187_ci_1 ));
    CascadeMux I__991 (
            .O(N__8995),
            .I(N__8991));
    InMux I__990 (
            .O(N__8994),
            .I(N__8988));
    InMux I__989 (
            .O(N__8991),
            .I(N__8985));
    LocalMux I__988 (
            .O(N__8988),
            .I(N__8981));
    LocalMux I__987 (
            .O(N__8985),
            .I(N__8978));
    InMux I__986 (
            .O(N__8984),
            .I(N__8975));
    Span4Mux_s1_h I__985 (
            .O(N__8981),
            .I(N__8972));
    Odrv4 I__984 (
            .O(N__8978),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__983 (
            .O(N__8975),
            .I(\uu0.l_countZ0Z_15 ));
    Odrv4 I__982 (
            .O(N__8972),
            .I(\uu0.l_countZ0Z_15 ));
    InMux I__981 (
            .O(N__8965),
            .I(N__8962));
    LocalMux I__980 (
            .O(N__8962),
            .I(\uu0.un4_l_count_12 ));
    CascadeMux I__979 (
            .O(N__8959),
            .I(N__8954));
    InMux I__978 (
            .O(N__8958),
            .I(N__8949));
    InMux I__977 (
            .O(N__8957),
            .I(N__8949));
    InMux I__976 (
            .O(N__8954),
            .I(N__8946));
    LocalMux I__975 (
            .O(N__8949),
            .I(\uu0.l_countZ0Z_17 ));
    LocalMux I__974 (
            .O(N__8946),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__973 (
            .O(N__8941),
            .I(N__8936));
    InMux I__972 (
            .O(N__8940),
            .I(N__8929));
    InMux I__971 (
            .O(N__8939),
            .I(N__8929));
    InMux I__970 (
            .O(N__8936),
            .I(N__8929));
    LocalMux I__969 (
            .O(N__8929),
            .I(N__8926));
    Odrv12 I__968 (
            .O(N__8926),
            .I(\uu0.un198_ci_2 ));
    CascadeMux I__967 (
            .O(N__8923),
            .I(N__8920));
    InMux I__966 (
            .O(N__8920),
            .I(N__8914));
    InMux I__965 (
            .O(N__8919),
            .I(N__8909));
    InMux I__964 (
            .O(N__8918),
            .I(N__8909));
    InMux I__963 (
            .O(N__8917),
            .I(N__8906));
    LocalMux I__962 (
            .O(N__8914),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__961 (
            .O(N__8909),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__960 (
            .O(N__8906),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__959 (
            .O(N__8899),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__958 (
            .O(N__8896),
            .I(N__8892));
    InMux I__957 (
            .O(N__8895),
            .I(N__8889));
    LocalMux I__956 (
            .O(N__8892),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__955 (
            .O(N__8889),
            .I(\uu0.l_countZ0Z_18 ));
    CascadeMux I__954 (
            .O(N__8884),
            .I(N__8878));
    CascadeMux I__953 (
            .O(N__8883),
            .I(N__8873));
    CascadeMux I__952 (
            .O(N__8882),
            .I(N__8870));
    InMux I__951 (
            .O(N__8881),
            .I(N__8863));
    InMux I__950 (
            .O(N__8878),
            .I(N__8856));
    InMux I__949 (
            .O(N__8877),
            .I(N__8856));
    InMux I__948 (
            .O(N__8876),
            .I(N__8856));
    InMux I__947 (
            .O(N__8873),
            .I(N__8847));
    InMux I__946 (
            .O(N__8870),
            .I(N__8847));
    InMux I__945 (
            .O(N__8869),
            .I(N__8847));
    InMux I__944 (
            .O(N__8868),
            .I(N__8847));
    InMux I__943 (
            .O(N__8867),
            .I(N__8842));
    InMux I__942 (
            .O(N__8866),
            .I(N__8842));
    LocalMux I__941 (
            .O(N__8863),
            .I(N__8835));
    LocalMux I__940 (
            .O(N__8856),
            .I(N__8835));
    LocalMux I__939 (
            .O(N__8847),
            .I(N__8835));
    LocalMux I__938 (
            .O(N__8842),
            .I(\uu0.un110_ci ));
    Odrv4 I__937 (
            .O(N__8835),
            .I(\uu0.un110_ci ));
    InMux I__936 (
            .O(N__8830),
            .I(N__8822));
    InMux I__935 (
            .O(N__8829),
            .I(N__8811));
    InMux I__934 (
            .O(N__8828),
            .I(N__8811));
    InMux I__933 (
            .O(N__8827),
            .I(N__8811));
    InMux I__932 (
            .O(N__8826),
            .I(N__8811));
    InMux I__931 (
            .O(N__8825),
            .I(N__8811));
    LocalMux I__930 (
            .O(N__8822),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__929 (
            .O(N__8811),
            .I(\uu0.l_countZ0Z_8 ));
    InMux I__928 (
            .O(N__8806),
            .I(N__8799));
    InMux I__927 (
            .O(N__8805),
            .I(N__8794));
    InMux I__926 (
            .O(N__8804),
            .I(N__8794));
    InMux I__925 (
            .O(N__8803),
            .I(N__8789));
    InMux I__924 (
            .O(N__8802),
            .I(N__8789));
    LocalMux I__923 (
            .O(N__8799),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__922 (
            .O(N__8794),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__921 (
            .O(N__8789),
            .I(\uu0.l_countZ0Z_9 ));
    CascadeMux I__920 (
            .O(N__8782),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__919 (
            .O(N__8779),
            .I(N__8770));
    InMux I__918 (
            .O(N__8778),
            .I(N__8770));
    InMux I__917 (
            .O(N__8777),
            .I(N__8770));
    LocalMux I__916 (
            .O(N__8770),
            .I(\uu2.l_countZ0Z_3 ));
    InMux I__915 (
            .O(N__8767),
            .I(N__8760));
    InMux I__914 (
            .O(N__8766),
            .I(N__8751));
    InMux I__913 (
            .O(N__8765),
            .I(N__8751));
    InMux I__912 (
            .O(N__8764),
            .I(N__8751));
    InMux I__911 (
            .O(N__8763),
            .I(N__8751));
    LocalMux I__910 (
            .O(N__8760),
            .I(N__8746));
    LocalMux I__909 (
            .O(N__8751),
            .I(N__8746));
    Odrv4 I__908 (
            .O(N__8746),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__907 (
            .O(N__8743),
            .I(N__8737));
    InMux I__906 (
            .O(N__8742),
            .I(N__8734));
    InMux I__905 (
            .O(N__8741),
            .I(N__8729));
    InMux I__904 (
            .O(N__8740),
            .I(N__8729));
    LocalMux I__903 (
            .O(N__8737),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__902 (
            .O(N__8734),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__901 (
            .O(N__8729),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__900 (
            .O(N__8722),
            .I(\uu0.un165_ci_0_cascade_ ));
    InMux I__899 (
            .O(N__8719),
            .I(N__8713));
    InMux I__898 (
            .O(N__8718),
            .I(N__8713));
    LocalMux I__897 (
            .O(N__8713),
            .I(\uu0.l_countZ0Z_13 ));
    CascadeMux I__896 (
            .O(N__8710),
            .I(N__8707));
    InMux I__895 (
            .O(N__8707),
            .I(N__8701));
    InMux I__894 (
            .O(N__8706),
            .I(N__8698));
    InMux I__893 (
            .O(N__8705),
            .I(N__8695));
    InMux I__892 (
            .O(N__8704),
            .I(N__8692));
    LocalMux I__891 (
            .O(N__8701),
            .I(N__8689));
    LocalMux I__890 (
            .O(N__8698),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__889 (
            .O(N__8695),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__888 (
            .O(N__8692),
            .I(\uu0.un154_ci_9 ));
    Odrv4 I__887 (
            .O(N__8689),
            .I(\uu0.un154_ci_9 ));
    CascadeMux I__886 (
            .O(N__8680),
            .I(\uu0.un110_ci_cascade_ ));
    InMux I__885 (
            .O(N__8677),
            .I(N__8668));
    InMux I__884 (
            .O(N__8676),
            .I(N__8668));
    InMux I__883 (
            .O(N__8675),
            .I(N__8668));
    LocalMux I__882 (
            .O(N__8668),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__881 (
            .O(N__8665),
            .I(N__8659));
    InMux I__880 (
            .O(N__8664),
            .I(N__8652));
    InMux I__879 (
            .O(N__8663),
            .I(N__8652));
    InMux I__878 (
            .O(N__8662),
            .I(N__8652));
    LocalMux I__877 (
            .O(N__8659),
            .I(N__8649));
    LocalMux I__876 (
            .O(N__8652),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__875 (
            .O(N__8649),
            .I(\uu0.l_countZ0Z_6 ));
    CascadeMux I__874 (
            .O(N__8644),
            .I(N__8639));
    InMux I__873 (
            .O(N__8643),
            .I(N__8636));
    InMux I__872 (
            .O(N__8642),
            .I(N__8631));
    InMux I__871 (
            .O(N__8639),
            .I(N__8631));
    LocalMux I__870 (
            .O(N__8636),
            .I(\uu2.l_countZ0Z_9 ));
    LocalMux I__869 (
            .O(N__8631),
            .I(\uu2.l_countZ0Z_9 ));
    CascadeMux I__868 (
            .O(N__8626),
            .I(N__8620));
    InMux I__867 (
            .O(N__8625),
            .I(N__8608));
    InMux I__866 (
            .O(N__8624),
            .I(N__8608));
    InMux I__865 (
            .O(N__8623),
            .I(N__8608));
    InMux I__864 (
            .O(N__8620),
            .I(N__8608));
    InMux I__863 (
            .O(N__8619),
            .I(N__8608));
    LocalMux I__862 (
            .O(N__8608),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__861 (
            .O(N__8605),
            .I(N__8598));
    InMux I__860 (
            .O(N__8604),
            .I(N__8598));
    InMux I__859 (
            .O(N__8603),
            .I(N__8595));
    LocalMux I__858 (
            .O(N__8598),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__857 (
            .O(N__8595),
            .I(\uu2.l_countZ0Z_5 ));
    CascadeMux I__856 (
            .O(N__8590),
            .I(N__8585));
    InMux I__855 (
            .O(N__8589),
            .I(N__8582));
    InMux I__854 (
            .O(N__8588),
            .I(N__8579));
    InMux I__853 (
            .O(N__8585),
            .I(N__8576));
    LocalMux I__852 (
            .O(N__8582),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__851 (
            .O(N__8579),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__850 (
            .O(N__8576),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__849 (
            .O(N__8569),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    InMux I__848 (
            .O(N__8566),
            .I(N__8563));
    LocalMux I__847 (
            .O(N__8563),
            .I(\uu2.un1_l_count_1_2_0 ));
    InMux I__846 (
            .O(N__8560),
            .I(N__8554));
    CascadeMux I__845 (
            .O(N__8559),
            .I(N__8551));
    InMux I__844 (
            .O(N__8558),
            .I(N__8548));
    InMux I__843 (
            .O(N__8557),
            .I(N__8545));
    LocalMux I__842 (
            .O(N__8554),
            .I(N__8542));
    InMux I__841 (
            .O(N__8551),
            .I(N__8539));
    LocalMux I__840 (
            .O(N__8548),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__839 (
            .O(N__8545),
            .I(\uu0.l_countZ0Z_14 ));
    Odrv4 I__838 (
            .O(N__8542),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__837 (
            .O(N__8539),
            .I(\uu0.l_countZ0Z_14 ));
    InMux I__836 (
            .O(N__8530),
            .I(N__8527));
    LocalMux I__835 (
            .O(N__8527),
            .I(\uu2.un1_l_count_2_2 ));
    InMux I__834 (
            .O(N__8524),
            .I(N__8521));
    LocalMux I__833 (
            .O(N__8521),
            .I(\uu2.un1_l_count_1_3 ));
    InMux I__832 (
            .O(N__8518),
            .I(N__8513));
    InMux I__831 (
            .O(N__8517),
            .I(N__8508));
    InMux I__830 (
            .O(N__8516),
            .I(N__8508));
    LocalMux I__829 (
            .O(N__8513),
            .I(N__8505));
    LocalMux I__828 (
            .O(N__8508),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__827 (
            .O(N__8505),
            .I(\uu2.un1_l_count_2_0 ));
    InMux I__826 (
            .O(N__8500),
            .I(N__8497));
    LocalMux I__825 (
            .O(N__8497),
            .I(vbuf_tx_data_2));
    InMux I__824 (
            .O(N__8494),
            .I(N__8491));
    LocalMux I__823 (
            .O(N__8491),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__822 (
            .O(N__8488),
            .I(N__8485));
    LocalMux I__821 (
            .O(N__8485),
            .I(vbuf_tx_data_3));
    InMux I__820 (
            .O(N__8482),
            .I(N__8479));
    LocalMux I__819 (
            .O(N__8479),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__818 (
            .O(N__8476),
            .I(N__8473));
    LocalMux I__817 (
            .O(N__8473),
            .I(vbuf_tx_data_4));
    InMux I__816 (
            .O(N__8470),
            .I(N__8467));
    LocalMux I__815 (
            .O(N__8467),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__814 (
            .O(N__8464),
            .I(N__8461));
    LocalMux I__813 (
            .O(N__8461),
            .I(vbuf_tx_data_5));
    InMux I__812 (
            .O(N__8458),
            .I(N__8455));
    LocalMux I__811 (
            .O(N__8455),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__810 (
            .O(N__8452),
            .I(\uu2.vbuf_count.un328_ci_3_cascade_ ));
    InMux I__809 (
            .O(N__8449),
            .I(N__8446));
    LocalMux I__808 (
            .O(N__8446),
            .I(\uu2.un350_ci ));
    CascadeMux I__807 (
            .O(N__8443),
            .I(\uu2.un350_ci_cascade_ ));
    InMux I__806 (
            .O(N__8440),
            .I(N__8437));
    LocalMux I__805 (
            .O(N__8437),
            .I(\uu2.r_data_wire_3 ));
    InMux I__804 (
            .O(N__8434),
            .I(N__8431));
    LocalMux I__803 (
            .O(N__8431),
            .I(\uu2.r_data_wire_4 ));
    InMux I__802 (
            .O(N__8428),
            .I(N__8425));
    LocalMux I__801 (
            .O(N__8425),
            .I(\uu2.r_data_wire_5 ));
    InMux I__800 (
            .O(N__8422),
            .I(N__8419));
    LocalMux I__799 (
            .O(N__8419),
            .I(\uu2.r_data_wire_6 ));
    InMux I__798 (
            .O(N__8416),
            .I(N__8413));
    LocalMux I__797 (
            .O(N__8413),
            .I(\uu2.r_data_wire_7 ));
    InMux I__796 (
            .O(N__8410),
            .I(N__8407));
    LocalMux I__795 (
            .O(N__8407),
            .I(vbuf_tx_data_0));
    InMux I__794 (
            .O(N__8404),
            .I(N__8401));
    LocalMux I__793 (
            .O(N__8401),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__792 (
            .O(N__8398),
            .I(N__8395));
    LocalMux I__791 (
            .O(N__8395),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__790 (
            .O(N__8392),
            .I(N__8389));
    LocalMux I__789 (
            .O(N__8389),
            .I(N__8386));
    Span12Mux_s1_h I__788 (
            .O(N__8386),
            .I(N__8383));
    Odrv12 I__787 (
            .O(N__8383),
            .I(o_serial_data_c));
    InMux I__786 (
            .O(N__8380),
            .I(N__8377));
    LocalMux I__785 (
            .O(N__8377),
            .I(vbuf_tx_data_1));
    InMux I__784 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__783 (
            .O(N__8371),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__782 (
            .O(N__8368),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__781 (
            .O(N__8365),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    CascadeMux I__780 (
            .O(N__8362),
            .I(N__8357));
    InMux I__779 (
            .O(N__8361),
            .I(N__8352));
    InMux I__778 (
            .O(N__8360),
            .I(N__8343));
    InMux I__777 (
            .O(N__8357),
            .I(N__8343));
    InMux I__776 (
            .O(N__8356),
            .I(N__8343));
    InMux I__775 (
            .O(N__8355),
            .I(N__8343));
    LocalMux I__774 (
            .O(N__8352),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__773 (
            .O(N__8343),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    InMux I__772 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__771 (
            .O(N__8335),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__770 (
            .O(N__8332),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__769 (
            .O(N__8329),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__768 (
            .O(N__8326),
            .I(N__8323));
    InMux I__767 (
            .O(N__8323),
            .I(N__8317));
    InMux I__766 (
            .O(N__8322),
            .I(N__8310));
    InMux I__765 (
            .O(N__8321),
            .I(N__8310));
    InMux I__764 (
            .O(N__8320),
            .I(N__8310));
    LocalMux I__763 (
            .O(N__8317),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__762 (
            .O(N__8310),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__761 (
            .O(N__8305),
            .I(N__8302));
    InMux I__760 (
            .O(N__8302),
            .I(N__8299));
    LocalMux I__759 (
            .O(N__8299),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__758 (
            .O(N__8296),
            .I(N__8285));
    InMux I__757 (
            .O(N__8295),
            .I(N__8285));
    InMux I__756 (
            .O(N__8294),
            .I(N__8285));
    InMux I__755 (
            .O(N__8293),
            .I(N__8282));
    InMux I__754 (
            .O(N__8292),
            .I(N__8279));
    LocalMux I__753 (
            .O(N__8285),
            .I(N__8276));
    LocalMux I__752 (
            .O(N__8282),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__751 (
            .O(N__8279),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    Odrv4 I__750 (
            .O(N__8276),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    InMux I__749 (
            .O(N__8269),
            .I(N__8266));
    LocalMux I__748 (
            .O(N__8266),
            .I(\uu2.r_data_wire_0 ));
    InMux I__747 (
            .O(N__8263),
            .I(N__8260));
    LocalMux I__746 (
            .O(N__8260),
            .I(\uu2.r_data_wire_1 ));
    InMux I__745 (
            .O(N__8257),
            .I(N__8254));
    LocalMux I__744 (
            .O(N__8254),
            .I(\uu2.r_data_wire_2 ));
    InMux I__743 (
            .O(N__8251),
            .I(N__8244));
    InMux I__742 (
            .O(N__8250),
            .I(N__8237));
    InMux I__741 (
            .O(N__8249),
            .I(N__8237));
    InMux I__740 (
            .O(N__8248),
            .I(N__8237));
    InMux I__739 (
            .O(N__8247),
            .I(N__8233));
    LocalMux I__738 (
            .O(N__8244),
            .I(N__8228));
    LocalMux I__737 (
            .O(N__8237),
            .I(N__8228));
    InMux I__736 (
            .O(N__8236),
            .I(N__8225));
    LocalMux I__735 (
            .O(N__8233),
            .I(N__8222));
    Odrv12 I__734 (
            .O(N__8228),
            .I(\uu0.l_precountZ0Z_0 ));
    LocalMux I__733 (
            .O(N__8225),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__732 (
            .O(N__8222),
            .I(\uu0.l_precountZ0Z_0 ));
    InMux I__731 (
            .O(N__8215),
            .I(N__8208));
    InMux I__730 (
            .O(N__8214),
            .I(N__8199));
    InMux I__729 (
            .O(N__8213),
            .I(N__8199));
    InMux I__728 (
            .O(N__8212),
            .I(N__8199));
    InMux I__727 (
            .O(N__8211),
            .I(N__8199));
    LocalMux I__726 (
            .O(N__8208),
            .I(\uu0.l_precountZ0Z_1 ));
    LocalMux I__725 (
            .O(N__8199),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__724 (
            .O(N__8194),
            .I(\buart.Z_rx.idle_0_cascade_ ));
    CascadeMux I__723 (
            .O(N__8191),
            .I(\buart.Z_rx.valid_0_cascade_ ));
    CascadeMux I__722 (
            .O(N__8188),
            .I(bu_rx_data_rdy_cascade_));
    CascadeMux I__721 (
            .O(N__8185),
            .I(\buart.Z_rx.N_27_0_i_cascade_ ));
    CascadeMux I__720 (
            .O(N__8182),
            .I(\uu0.un143_ci_0_cascade_ ));
    CascadeMux I__719 (
            .O(N__8179),
            .I(\uu0.un4_l_count_11_cascade_ ));
    InMux I__718 (
            .O(N__8176),
            .I(N__8173));
    LocalMux I__717 (
            .O(N__8173),
            .I(\uu0.un4_l_count_18 ));
    CascadeMux I__716 (
            .O(N__8170),
            .I(\uu0.un4_l_count_16_cascade_ ));
    CascadeMux I__715 (
            .O(N__8167),
            .I(N__8162));
    CascadeMux I__714 (
            .O(N__8166),
            .I(N__8159));
    InMux I__713 (
            .O(N__8165),
            .I(N__8152));
    InMux I__712 (
            .O(N__8162),
            .I(N__8152));
    InMux I__711 (
            .O(N__8159),
            .I(N__8152));
    LocalMux I__710 (
            .O(N__8152),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__709 (
            .O(N__8149),
            .I(N__8146));
    InMux I__708 (
            .O(N__8146),
            .I(N__8134));
    InMux I__707 (
            .O(N__8145),
            .I(N__8134));
    InMux I__706 (
            .O(N__8144),
            .I(N__8134));
    InMux I__705 (
            .O(N__8143),
            .I(N__8134));
    LocalMux I__704 (
            .O(N__8134),
            .I(\uu0.l_precountZ0Z_2 ));
    CascadeMux I__703 (
            .O(N__8131),
            .I(N__8127));
    InMux I__702 (
            .O(N__8130),
            .I(N__8121));
    InMux I__701 (
            .O(N__8127),
            .I(N__8121));
    InMux I__700 (
            .O(N__8126),
            .I(N__8118));
    LocalMux I__699 (
            .O(N__8121),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__698 (
            .O(N__8118),
            .I(\uu0.l_countZ0Z_11 ));
    InMux I__697 (
            .O(N__8113),
            .I(N__8110));
    LocalMux I__696 (
            .O(N__8110),
            .I(\uu0.un4_l_count_13 ));
    CascadeMux I__695 (
            .O(N__8107),
            .I(\uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__694 (
            .O(N__8104),
            .I(\uu0.un154_ci_9_cascade_ ));
    InMux I__693 (
            .O(N__8101),
            .I(N__8089));
    InMux I__692 (
            .O(N__8100),
            .I(N__8089));
    InMux I__691 (
            .O(N__8099),
            .I(N__8089));
    InMux I__690 (
            .O(N__8098),
            .I(N__8089));
    LocalMux I__689 (
            .O(N__8089),
            .I(\uu0.l_countZ0Z_10 ));
    IoInMux I__688 (
            .O(N__8086),
            .I(N__8083));
    LocalMux I__687 (
            .O(N__8083),
            .I(N__8080));
    Span12Mux_s9_v I__686 (
            .O(N__8080),
            .I(N__8077));
    Odrv12 I__685 (
            .O(N__8077),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__684 (
            .O(N__8074),
            .I(N__8071));
    LocalMux I__683 (
            .O(N__8071),
            .I(N__8068));
    IoSpan4Mux I__682 (
            .O(N__8068),
            .I(N__8065));
    Odrv4 I__681 (
            .O(N__8065),
            .I(clk_in_c));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__22339));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__22342));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__22346));
    INV \INVuu2.bitmap_215C  (
            .O(\INVuu2.bitmap_215C_net ),
            .I(N__22321));
    INV \INVuu2.w_addr_displaying_7C  (
            .O(\INVuu2.w_addr_displaying_7C_net ),
            .I(N__22338));
    INV \INVuu2.w_addr_displaying_ness_6C  (
            .O(\INVuu2.w_addr_displaying_ness_6C_net ),
            .I(N__22341));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__22320));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__22325));
    INV \INVuu2.bitmap_40C  (
            .O(\INVuu2.bitmap_40C_net ),
            .I(N__22332));
    INV \INVuu2.w_addr_displaying_fast_8C  (
            .O(\INVuu2.w_addr_displaying_fast_8C_net ),
            .I(N__22337));
    INV \INVuu2.bitmap_197C  (
            .O(\INVuu2.bitmap_197C_net ),
            .I(N__22315));
    INV \INVuu2.w_addr_displaying_1_rep1_nesrC  (
            .O(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .I(N__22323));
    INV \INVuu2.w_addr_user_2C  (
            .O(\INVuu2.w_addr_user_2C_net ),
            .I(N__22327));
    INV \INVuu2.w_addr_displaying_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .I(N__22331));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__22348));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__8086),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__9433),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__9259),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__12723),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.l_count_8_LC_1_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_1_6_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_1_6_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__8588),
            .in2(_gnd_net_),
            .in3(N__8449),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22328),
            .ce(),
            .sr(N__20953));
    defparam \uu2.l_count_1_LC_1_6_3 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_1_6_3 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_1_6_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_1_LC_1_6_3  (
            .in0(N__10338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10372),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22328),
            .ce(),
            .sr(N__20953));
    defparam \uu2.l_count_0_LC_1_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_1_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10337),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22328),
            .ce(),
            .sr(N__20953));
    defparam \uu0.l_precount_0_LC_1_6_6 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_1_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8236),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22328),
            .ce(),
            .sr(N__20953));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_7_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_7_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_7_7  (
            .in0(N__8704),
            .in1(N__8557),
            .in2(_gnd_net_),
            .in3(N__8743),
            .lcout(\uu0.un187_ci_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI04591_10_LC_1_8_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI04591_10_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI04591_10_LC_1_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_count_RNI04591_10_LC_1_8_0  (
            .in0(N__8098),
            .in1(N__8825),
            .in2(N__8559),
            .in3(N__9169),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2GS72_4_LC_1_8_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_8_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNI2GS72_4_LC_1_8_1  (
            .in0(N__8247),
            .in1(N__8740),
            .in2(N__8107),
            .in3(N__9052),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_10_LC_1_8_2 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_8_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_10_LC_1_8_2  (
            .in0(N__8101),
            .in1(N__8806),
            .in2(N__8884),
            .in3(N__8828),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(N__9074),
            .sr(N__20949));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_8_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_8_3  (
            .in0(N__8826),
            .in1(N__8804),
            .in2(N__8131),
            .in3(N__8099),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_1_8_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_8_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_1_8_4  (
            .in0(N__8741),
            .in1(N__8558),
            .in2(N__8104),
            .in3(N__8881),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(N__9074),
            .sr(N__20949));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_8_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_8_5  (
            .in0(N__8827),
            .in1(N__8805),
            .in2(_gnd_net_),
            .in3(N__8100),
            .lcout(),
            .ltout(\uu0.un143_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_11_LC_1_8_6 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_1_8_6 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_11_LC_1_8_6  (
            .in0(N__8877),
            .in1(N__8130),
            .in2(N__8182),
            .in3(N__9323),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(N__9074),
            .sr(N__20949));
    defparam \uu0.l_count_8_LC_1_8_7 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_8_LC_1_8_7  (
            .in0(N__8829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(N__9074),
            .sr(N__20949));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_0 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_9_0  (
            .in0(N__8211),
            .in1(N__9035),
            .in2(N__8166),
            .in3(N__9121),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI96A32_18_LC_1_9_1  (
            .in0(N__8665),
            .in1(N__8895),
            .in2(N__8179),
            .in3(N__8994),
            .lcout(),
            .ltout(\uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_11_LC_1_9_2  (
            .in0(N__8113),
            .in1(N__8176),
            .in2(N__8170),
            .in3(N__8965),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_2_LC_1_9_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_9_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu0.l_precount_2_LC_1_9_4  (
            .in0(N__8213),
            .in1(N__8145),
            .in2(_gnd_net_),
            .in3(N__8249),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(N__20951));
    defparam \uu0.l_precount_3_LC_1_9_5 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_9_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_9_5  (
            .in0(N__8250),
            .in1(N__8165),
            .in2(N__8149),
            .in3(N__8214),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(N__20951));
    defparam \uu0.delay_line_0_LC_1_9_6 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_9_6  (
            .in0(N__8212),
            .in1(N__8144),
            .in2(N__8167),
            .in3(N__8248),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(N__20951));
    defparam \uu0.l_count_RNI2CNU_11_LC_1_9_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_9_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNI2CNU_11_LC_1_9_7  (
            .in0(N__8143),
            .in1(N__8126),
            .in2(N__9150),
            .in3(N__8917),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_1_LC_1_10_0 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9349),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22300),
            .ce(),
            .sr(N__20952));
    defparam \uu0.l_precount_1_LC_1_10_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_precount_1_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__8251),
            .in2(_gnd_net_),
            .in3(N__8215),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22300),
            .ce(),
            .sr(N__20952));
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_11_0  (
            .in0(N__8322),
            .in1(N__9401),
            .in2(N__8362),
            .in3(N__8295),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__8355),
            .in2(_gnd_net_),
            .in3(N__8320),
            .lcout(),
            .ltout(\buart.Z_rx.idle_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_11_2  (
            .in0(N__9454),
            .in1(N__9399),
            .in2(N__8194),
            .in3(N__8296),
            .lcout(\buart.Z_rx.idle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__8321),
            .in2(_gnd_net_),
            .in3(N__9453),
            .lcout(),
            .ltout(\buart.Z_rx.valid_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_11_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_11_4  (
            .in0(N__8356),
            .in1(N__9400),
            .in2(N__8191),
            .in3(N__8294),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_1_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_1_11_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8188),
            .in3(N__13784),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(\buart.Z_rx.N_27_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_1_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_11_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_11_6 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_1_11_6  (
            .in0(N__8360),
            .in1(N__8338),
            .in2(N__8185),
            .in3(N__13759),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22291),
            .ce(N__9768),
            .sr(N__20956));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_12_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_12_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__8292),
            .in2(_gnd_net_),
            .in3(N__8368),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_12_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9409),
            .in3(N__8365),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_12_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__8361),
            .in2(_gnd_net_),
            .in3(N__8332),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_1_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_12_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_12_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_1_12_4  (
            .in0(N__9373),
            .in1(N__13757),
            .in2(N__8326),
            .in3(N__8329),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__9766),
            .sr(N__20959));
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .LUT_INIT=16'b0001010010111110;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_1_13_4  (
            .in0(N__9379),
            .in1(N__8293),
            .in2(N__8305),
            .in3(N__13760),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22277),
            .ce(N__9769),
            .sr(N__20961));
    defparam \uu2.r_data_reg_0_LC_2_1_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_0_LC_2_1_0  (
            .in0(N__8269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_1_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_1_LC_2_1_1  (
            .in0(N__8263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_1_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_2_LC_2_1_2  (
            .in0(N__8257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_1_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_3_LC_2_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8440),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_1_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8434),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_1_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8428),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_1_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8422),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_1_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_7_LC_2_1_7  (
            .in0(N__8416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_2_0  (
            .in0(N__21708),
            .in1(N__8374),
            .in2(_gnd_net_),
            .in3(N__8410),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__8404),
            .in2(_gnd_net_),
            .in3(N__21706),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_2_2  (
            .in0(N__21707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8398),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_2_3  (
            .in0(N__8494),
            .in1(N__21709),
            .in2(_gnd_net_),
            .in3(N__8380),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_2_4  (
            .in0(N__21710),
            .in1(N__8482),
            .in2(_gnd_net_),
            .in3(N__8500),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_2_5  (
            .in0(N__8488),
            .in1(N__8470),
            .in2(_gnd_net_),
            .in3(N__21711),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_2_6  (
            .in0(N__21712),
            .in1(N__8458),
            .in2(_gnd_net_),
            .in3(N__8476),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_2_7  (
            .in0(N__10444),
            .in1(N__21713),
            .in2(_gnd_net_),
            .in3(N__8464),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(N__21621),
            .sr(N__20964));
    defparam \uu0.sec_clk_LC_2_4_2 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_2_4_2 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_2_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__13546),
            .in2(_gnd_net_),
            .in3(N__9336),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22335),
            .ce(),
            .sr(N__20962));
    defparam \uu2.vram_rd_clk_LC_2_4_6 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_2_4_6 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_2_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(N__14347),
            .in2(_gnd_net_),
            .in3(N__8518),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22335),
            .ce(),
            .sr(N__20962));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_0 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__8623),
            .in2(_gnd_net_),
            .in3(N__8604),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(\uu2.vbuf_count.un328_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1  (
            .in0(N__10005),
            .in1(N__10070),
            .in2(N__8452),
            .in3(N__10023),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_2_5_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uu2.l_count_9_LC_2_5_2  (
            .in0(N__8517),
            .in1(N__8643),
            .in2(N__8443),
            .in3(N__8589),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__20960));
    defparam \uu2.l_count_4_LC_2_5_3 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_2_5_3 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_2_5_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu2.l_count_4_LC_2_5_3  (
            .in0(N__8624),
            .in1(N__10025),
            .in2(_gnd_net_),
            .in3(N__8516),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__20960));
    defparam \uu2.l_count_5_LC_2_5_4 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_2_5_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_5_LC_2_5_4  (
            .in0(N__10026),
            .in1(N__8625),
            .in2(_gnd_net_),
            .in3(N__8605),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__20960));
    defparam \uu2.l_count_6_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_2_5_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_2_5_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.l_count_6_LC_2_5_5  (
            .in0(N__10044),
            .in1(N__10071),
            .in2(_gnd_net_),
            .in3(N__10024),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__20960));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6  (
            .in0(N__10068),
            .in1(N__8619),
            .in2(N__8644),
            .in3(N__10331),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_2_5_7  (
            .in0(N__10332),
            .in1(N__8642),
            .in2(N__8626),
            .in3(N__10069),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_2_6_0  (
            .in0(N__8603),
            .in1(N__10006),
            .in2(N__8590),
            .in3(N__8777),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_2_6_1  (
            .in0(N__10365),
            .in1(N__8763),
            .in2(N__8569),
            .in3(N__8566),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2  (
            .in0(N__8984),
            .in1(N__8560),
            .in2(N__8710),
            .in3(N__8742),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_2_6_3  (
            .in0(N__8530),
            .in1(N__8765),
            .in2(N__10374),
            .in3(N__8524),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_3_LC_2_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_2_6_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uu2.l_count_3_LC_2_6_4  (
            .in0(N__10306),
            .in1(N__8767),
            .in2(N__8782),
            .in3(N__8779),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(N__20958));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6  (
            .in0(N__8764),
            .in1(N__8778),
            .in2(N__10373),
            .in3(N__10333),
            .lcout(\uu2.un306_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_2_6_7 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_2_6_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_2_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__10305),
            .in2(_gnd_net_),
            .in3(N__8766),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(N__20958));
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__8718),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_7_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_7_1  (
            .in0(N__8663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9020),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__8705),
            .in2(_gnd_net_),
            .in3(N__8676),
            .lcout(),
            .ltout(\uu0.un165_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_13_LC_2_7_3 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_2_7_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_2_7_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_13_LC_2_7_3  (
            .in0(N__8719),
            .in1(N__8866),
            .in2(N__8722),
            .in3(N__9331),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22317),
            .ce(N__9076),
            .sr(N__20954));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_7_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_7_4  (
            .in0(N__9099),
            .in1(N__8662),
            .in2(N__9022),
            .in3(N__9217),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_12_LC_2_7_5 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_2_7_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_2_7_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_12_LC_2_7_5  (
            .in0(N__8677),
            .in1(N__8706),
            .in2(N__8680),
            .in3(N__9330),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22317),
            .ce(N__9076),
            .sr(N__20954));
    defparam \uu0.l_count_6_LC_2_7_6 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_2_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_2_7_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_6_LC_2_7_6  (
            .in0(N__9021),
            .in1(N__9337),
            .in2(N__9103),
            .in3(N__8664),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22317),
            .ce(N__9076),
            .sr(N__20954));
    defparam \uu0.l_count_15_LC_2_7_7 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_2_7_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_15_LC_2_7_7  (
            .in0(N__9004),
            .in1(N__8867),
            .in2(N__8995),
            .in3(N__9332),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22317),
            .ce(N__9076),
            .sr(N__20954));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_8_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_8_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_8_0  (
            .in0(N__8802),
            .in1(N__9215),
            .in2(N__8959),
            .in3(N__9191),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_2_8_1 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_2_8_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_2_8_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_16_LC_2_8_1  (
            .in0(N__8939),
            .in1(N__8869),
            .in2(N__8923),
            .in3(N__9324),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.l_count_17_LC_2_8_2 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_8_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_8_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_17_LC_2_8_2  (
            .in0(N__8919),
            .in1(N__8940),
            .in2(N__8882),
            .in3(N__8958),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_8_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_8_3  (
            .in0(N__8957),
            .in1(N__8868),
            .in2(N__8941),
            .in3(N__8918),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_8_4 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_8_4 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uu0.l_count_18_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__9321),
            .in2(N__8899),
            .in3(N__8896),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.l_count_3_LC_2_8_5 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_2_8_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_3_LC_2_8_5  (
            .in0(N__9192),
            .in1(N__9202),
            .in2(N__9178),
            .in3(N__9326),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.l_count_9_LC_2_8_6 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_2_8_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_2_8_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu0.l_count_9_LC_2_8_6  (
            .in0(N__8803),
            .in1(_gnd_net_),
            .in2(N__8883),
            .in3(N__8830),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.l_count_7_LC_2_8_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_2_8_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_2_8_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_7_LC_2_8_7  (
            .in0(N__9216),
            .in1(N__9098),
            .in2(N__9226),
            .in3(N__9325),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22309),
            .ce(N__9075),
            .sr(N__20950));
    defparam \uu0.l_count_0_LC_2_9_0 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_2_9_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_2_9_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_2_9_0  (
            .in0(N__9148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9322),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(N__9073),
            .sr(N__20955));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_9_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_9_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_9_1  (
            .in0(N__9123),
            .in1(N__9147),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.un44_ci ),
            .ltout(\uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_2_9_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_2_9_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_2_9_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu0.l_count_2_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9196),
            .in3(N__9171),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(N__9073),
            .sr(N__20955));
    defparam \uu0.l_count_1_LC_2_9_3 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_2_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_2_9_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \uu0.l_count_1_LC_2_9_3  (
            .in0(N__9124),
            .in1(N__9149),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(N__9073),
            .sr(N__20955));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_9_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_9_4  (
            .in0(N__9193),
            .in1(N__9170),
            .in2(N__9151),
            .in3(N__9122),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_4_LC_2_9_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_2_9_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_2_9_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uu0.l_count_4_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__9320),
            .in2(N__9106),
            .in3(N__9054),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(N__9073),
            .sr(N__20955));
    defparam \uu0.l_count_5_LC_2_9_6 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_2_9_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_2_9_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu0.l_count_5_LC_2_9_6  (
            .in0(N__9037),
            .in1(_gnd_net_),
            .in2(N__9058),
            .in3(N__9097),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(N__9073),
            .sr(N__20955));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__9053),
            .in2(_gnd_net_),
            .in3(N__9036),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_0 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_2_10_0  (
            .in0(N__13748),
            .in1(N__9378),
            .in2(N__9421),
            .in3(N__9405),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22292),
            .ce(N__9767),
            .sr(N__20957));
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_2_10_1  (
            .in0(N__9377),
            .in1(N__13749),
            .in2(N__10838),
            .in3(N__9461),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22292),
            .ce(N__9767),
            .sr(N__20957));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_10_4 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__9568),
            .in2(_gnd_net_),
            .in3(N__9587),
            .lcout(\resetGen.un241_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_2_10_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_2_10_5  (
            .in0(N__9494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9549),
            .lcout(\resetGen.reset_count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_2_10_6  (
            .in0(N__9355),
            .in1(N__9348),
            .in2(_gnd_net_),
            .in3(N__9306),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7  (
            .in0(N__15976),
            .in1(N__11149),
            .in2(_gnd_net_),
            .in3(N__21868),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_2_11_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_2_11_0 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_2_11_0  (
            .in0(N__11833),
            .in1(N__9537),
            .in2(N__9574),
            .in3(N__9589),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_2_11_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_2_11_1 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_2_11_1  (
            .in0(N__9534),
            .in1(N__9570),
            .in2(_gnd_net_),
            .in3(N__11832),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_2_11_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_2_11_2 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \resetGen.reset_count_4_LC_2_11_2  (
            .in0(N__11836),
            .in1(N__9510),
            .in2(N__9538),
            .in3(N__9232),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_3 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_3  (
            .in0(N__9588),
            .in1(N__9569),
            .in2(_gnd_net_),
            .in3(N__9495),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_2_11_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_2_11_4 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_3_LC_2_11_4  (
            .in0(N__11835),
            .in1(N__9536),
            .in2(N__9553),
            .in3(N__9550),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_2_11_5 .C_ON=1'b0;
    defparam \resetGen.rst_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_2_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_2_11_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_2_11_6 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \resetGen.reset_count_2_LC_2_11_6  (
            .in0(N__11834),
            .in1(N__9535),
            .in2(N__9499),
            .in3(N__9511),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_11_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__14797),
            .in2(_gnd_net_),
            .in3(N__21034),
            .lcout(\Lab_UT.didp.regrce2.LdAStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_0  (
            .in0(N__9735),
            .in1(N__9716),
            .in2(_gnd_net_),
            .in3(N__13752),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_1  (
            .in0(N__9672),
            .in1(N__9656),
            .in2(N__9606),
            .in3(N__9734),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__9695),
            .in2(N__9481),
            .in3(N__9712),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__9478),
            .in2(N__9469),
            .in3(N__9465),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4  (
            .in0(N__9682),
            .in1(N__9696),
            .in2(N__13764),
            .in3(N__9628),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_5  (
            .in0(N__13751),
            .in1(_gnd_net_),
            .in2(N__9720),
            .in3(_gnd_net_),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_6  (
            .in0(N__9657),
            .in1(N__9629),
            .in2(N__9643),
            .in3(N__13753),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7  (
            .in0(N__13750),
            .in1(N__13785),
            .in2(N__9631),
            .in3(N__18040),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__9736),
            .in2(N__9721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__9697),
            .in2(_gnd_net_),
            .in3(N__9676),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2  (
            .in0(N__13765),
            .in1(N__9673),
            .in2(_gnd_net_),
            .in3(N__9661),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__22273),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__9658),
            .in2(_gnd_net_),
            .in3(N__9634),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4  (
            .in0(N__9630),
            .in1(N__13758),
            .in2(N__9607),
            .in3(N__9610),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_1_0  (
            .in0(N__9927),
            .in1(N__9896),
            .in2(N__9831),
            .in3(N__10260),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__10228),
            .sr(N__20948));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_1 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(N__9845),
            .in2(_gnd_net_),
            .in3(N__9799),
            .lcout(),
            .ltout(\uu2.vbuf_raddr.un448_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_1_2  (
            .in0(N__10165),
            .in1(N__9861),
            .in2(N__9868),
            .in3(N__9783),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__10228),
            .sr(N__20948));
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_1_3  (
            .in0(N__9784),
            .in1(N__9846),
            .in2(N__10171),
            .in3(N__9800),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__10228),
            .sr(N__20948));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4  (
            .in0(N__9926),
            .in1(N__9895),
            .in2(N__9830),
            .in3(N__10259),
            .lcout(\uu2.un404_ci_0 ),
            .ltout(\uu2.un404_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_1_5  (
            .in0(N__10205),
            .in1(N__10117),
            .in2(N__9808),
            .in3(N__9801),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__10228),
            .sr(N__20948));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_6 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_6  (
            .in0(_gnd_net_),
            .in1(N__10103),
            .in2(_gnd_net_),
            .in3(N__10204),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7  (
            .in0(N__13228),
            .in1(N__13108),
            .in2(N__11896),
            .in3(N__13177),
            .lcout(\uu2.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0  (
            .in0(N__21911),
            .in1(N__12810),
            .in2(N__10537),
            .in3(N__10741),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1  (
            .in0(N__9973),
            .in1(N__10699),
            .in2(_gnd_net_),
            .in3(N__21910),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2  (
            .in0(N__10512),
            .in1(N__10529),
            .in2(_gnd_net_),
            .in3(N__12808),
            .lcout(\uu2.N_34 ),
            .ltout(\uu2.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3  (
            .in0(N__10894),
            .in1(N__21913),
            .in2(N__9967),
            .in3(N__10566),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4  (
            .in0(N__10567),
            .in1(N__9946),
            .in2(N__21919),
            .in3(N__10783),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5  (
            .in0(N__9945),
            .in1(N__10762),
            .in2(_gnd_net_),
            .in3(N__21909),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6  (
            .in0(N__10513),
            .in1(N__12809),
            .in2(N__10536),
            .in3(N__11148),
            .lcout(\uu2.N_31 ),
            .ltout(\uu2.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(N__21912),
            .in2(N__9937),
            .in3(N__11713),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_2_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_4_3_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_2_LC_4_3_0  (
            .in0(N__10140),
            .in1(N__9922),
            .in2(N__9900),
            .in3(N__10255),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(),
            .sr(N__20941));
    defparam \uu2.r_addr_1_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_4_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_1_LC_4_3_1  (
            .in0(N__10254),
            .in1(N__9891),
            .in2(_gnd_net_),
            .in3(N__10138),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(),
            .sr(N__20941));
    defparam \uu2.r_addr_0_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.r_addr_0_LC_4_3_2  (
            .in0(N__10137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10253),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(),
            .sr(N__20941));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__10136),
            .in2(_gnd_net_),
            .in3(N__21036),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_4_LC_4_3_7 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_3_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_4_3_7  (
            .in0(N__10197),
            .in1(N__10167),
            .in2(_gnd_net_),
            .in3(N__10139),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(),
            .sr(N__20941));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__11512),
            .in2(_gnd_net_),
            .in3(N__21885),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__10642),
            .in2(_gnd_net_),
            .in3(N__10635),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_5_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_4_5_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_4_5_0  (
            .in0(N__10206),
            .in1(N__10166),
            .in2(N__10102),
            .in3(N__10141),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__20934));
    defparam \uu2.l_count_7_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_4_5_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_4_5_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.l_count_7_LC_4_5_1  (
            .in0(N__10075),
            .in1(N__10001),
            .in2(N__10051),
            .in3(N__10033),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__20934));
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_4_5_2  (
            .in0(N__11206),
            .in1(_gnd_net_),
            .in2(N__12133),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__20934));
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__12129),
            .in2(_gnd_net_),
            .in3(N__11205),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__20934));
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__14704),
            .in2(_gnd_net_),
            .in3(N__21033),
            .lcout(\Lab_UT.didp.regrce3.LdAMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_6_2 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__10375),
            .in2(_gnd_net_),
            .in3(N__10339),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_6_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_6_5  (
            .in0(N__17650),
            .in1(N__17688),
            .in2(_gnd_net_),
            .in3(N__14258),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_4_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_4_6_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_4_6_6  (
            .in0(N__17689),
            .in1(N__17312),
            .in2(N__10294),
            .in3(N__17763),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22310),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_4_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_4_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_3_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20521),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22302),
            .ce(N__10291),
            .sr(N__20932));
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_4_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_4_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_0_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14259),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22302),
            .ce(N__10291),
            .sr(N__20932));
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_4_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_4_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_2_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20338),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22302),
            .ce(N__10291),
            .sr(N__20932));
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_4_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_1_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20154),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22293),
            .ce(N__10290),
            .sr(N__20931));
    defparam \Lab_UT.alarmchar_latch_6_LC_4_9_0 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_6_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_6_LC_4_9_0 .LUT_INIT=16'b0000000011011010;
    LogicCell40 \Lab_UT.alarmchar_latch_6_LC_4_9_0  (
            .in0(N__11414),
            .in1(N__10270),
            .in2(N__11358),
            .in3(N__10501),
            .lcout(G_184),
            .ltout(G_184_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_4_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_4_9_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_4_9_1  (
            .in0(N__18364),
            .in1(_gnd_net_),
            .in2(N__10264),
            .in3(N__11575),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22286),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_4_9_2 .C_ON=1'b0;
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_4_9_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \Lab_UT.un1_idle_1_0_iclk_LC_4_9_2  (
            .in0(N__11348),
            .in1(N__11411),
            .in2(_gnd_net_),
            .in3(N__21035),
            .lcout(),
            .ltout(\Lab_UT.un1_idle_1_0_iclkZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_3 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \Lab_UT.alarmchar_latch_3_LC_4_9_3  (
            .in0(N__10820),
            .in1(N__10915),
            .in2(N__10396),
            .in3(N__10479),
            .lcout(G_188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m59_LC_4_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m59_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m59_LC_4_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.m59_LC_4_9_5  (
            .in0(N__11410),
            .in1(N__12722),
            .in2(_gnd_net_),
            .in3(N__11347),
            .lcout(\Lab_UT.alarmstate_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_4_9_6  (
            .in0(N__11574),
            .in1(N__18363),
            .in2(_gnd_net_),
            .in3(N__10467),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_4_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_4_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_4_9_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_4_9_7  (
            .in0(N__13638),
            .in1(N__11599),
            .in2(N__10393),
            .in3(N__11746),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22286),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_4_10_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_4_10_0  (
            .in0(N__11407),
            .in1(N__21023),
            .in2(_gnd_net_),
            .in3(N__11343),
            .lcout(G_180),
            .ltout(G_180_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_4_10_1 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_1_LC_4_10_1  (
            .in0(N__11346),
            .in1(N__10500),
            .in2(N__10390),
            .in3(N__10951),
            .lcout(G_181),
            .ltout(G_181_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_4_10_2 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_0__m3_LC_4_10_2  (
            .in0(N__10942),
            .in1(N__12397),
            .in2(N__10387),
            .in3(N__11415),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_4_10_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_0_LC_4_10_3  (
            .in0(N__10384),
            .in1(N__11408),
            .in2(N__10378),
            .in3(N__10498),
            .lcout(G_179),
            .ltout(G_179_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_10_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.un1_armed_2_0_iso_i_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10504),
            .in3(N__11344),
            .lcout(\Lab_UT.un1_armed_2_0_iso_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_4_10_5 .C_ON=1'b0;
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_4_10_5 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \Lab_UT.un1_idle_5_0_iclk_LC_4_10_5  (
            .in0(N__11345),
            .in1(N__11409),
            .in2(_gnd_net_),
            .in3(N__10499),
            .lcout(),
            .ltout(\Lab_UT.un1_idle_5_0_iclkZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_1_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_1_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_1_LC_4_10_6 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \Lab_UT.alarmchar_latch_1_LC_4_10_6  (
            .in0(N__10468),
            .in1(N__10819),
            .in2(N__10483),
            .in3(N__10480),
            .lcout(G_185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_4_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_4_11_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20326),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22274),
            .ce(N__15481),
            .sr(N__20963));
    defparam \buart.Z_rx.shifter_0_LC_4_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_4_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_4_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20110),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22271),
            .ce(N__15480),
            .sr(N__20965));
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_5_1_0  (
            .in0(N__21697),
            .in1(N__10423),
            .in2(_gnd_net_),
            .in3(N__10456),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(N__21622),
            .sr(N__20971));
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__21696),
            .in2(_gnd_net_),
            .in3(N__10432),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(N__21622),
            .sr(N__20971));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2  (
            .in0(N__15871),
            .in1(N__21867),
            .in2(_gnd_net_),
            .in3(N__13338),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3  (
            .in0(N__13516),
            .in1(N__13498),
            .in2(_gnd_net_),
            .in3(N__21021),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4  (
            .in0(N__21791),
            .in1(N__20682),
            .in2(_gnd_net_),
            .in3(N__13176),
            .lcout(\uu2.w_addr_displaying_RNI03P31Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5  (
            .in0(N__16153),
            .in1(N__11488),
            .in2(_gnd_net_),
            .in3(N__10795),
            .lcout(\uu2.un28_w_addr_user_i ),
            .ltout(\uu2.un28_w_addr_user_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_user_RNID65PE_4_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10540),
            .in3(N__15822),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \uu2.w_addr_user_RNI43E87_4_LC_5_1_7  (
            .in0(N__16152),
            .in1(N__21020),
            .in2(_gnd_net_),
            .in3(N__10794),
            .lcout(\uu2.w_addr_user_RNI43E87Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_5_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_5_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIKIPH1_8_LC_5_2_0  (
            .in0(N__20684),
            .in1(N__21782),
            .in2(N__16136),
            .in3(N__13342),
            .lcout(\uu2.un51_w_data_displaying_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_5_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_5_2_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__11119),
            .in2(_gnd_net_),
            .in3(N__20683),
            .lcout(),
            .ltout(\uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_5_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_5_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIASLS1_8_LC_5_2_2  (
            .in0(N__21781),
            .in1(N__16126),
            .in2(N__10516),
            .in3(N__13341),
            .lcout(\uu2.w_data_displaying_2_i_a2_i_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_2_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_5_2_3  (
            .in0(N__16127),
            .in1(N__20687),
            .in2(N__21792),
            .in3(N__11124),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__13253),
            .sr(N__20895));
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_5_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_5_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_5_2_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_3_LC_5_2_4  (
            .in0(N__20685),
            .in1(N__21784),
            .in2(N__11135),
            .in3(N__11943),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__13253),
            .sr(N__20895));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_5_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_5_2_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_LC_5_2_5  (
            .in0(N__21783),
            .in1(N__20686),
            .in2(N__16468),
            .in3(N__11120),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__13253),
            .sr(N__20895));
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_5_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_5_2_6 .LUT_INIT=16'b1100110001001000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_5_2_6  (
            .in0(N__21780),
            .in1(N__12001),
            .in2(N__16135),
            .in3(N__11029),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_5_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_5_2_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_RNI0FGN6_4_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__10585),
            .in2(N__10579),
            .in3(N__11059),
            .lcout(\uu2.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0  (
            .in0(N__10648),
            .in1(N__10552),
            .in2(_gnd_net_),
            .in3(N__11014),
            .lcout(),
            .ltout(\uu2.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1  (
            .in0(N__10576),
            .in1(N__10546),
            .in2(N__10570),
            .in3(N__12013),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2  (
            .in0(N__16457),
            .in1(N__13339),
            .in2(_gnd_net_),
            .in3(N__12104),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNICM7R_180_LC_5_3_3  (
            .in0(N__16780),
            .in1(N__12190),
            .in2(_gnd_net_),
            .in3(N__11947),
            .lcout(),
            .ltout(\uu2.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4  (
            .in0(N__16458),
            .in1(N__16332),
            .in2(N__10558),
            .in3(N__12166),
            .lcout(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ),
            .ltout(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5  (
            .in0(N__11049),
            .in1(N__10665),
            .in2(N__10555),
            .in3(N__16731),
            .lcout(\uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6  (
            .in0(N__13340),
            .in1(N__11035),
            .in2(_gnd_net_),
            .in3(N__16333),
            .lcout(\uu2.bitmap_pmux_u_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .LUT_INIT=16'b1101111110001111;
    LogicCell40 \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7  (
            .in0(N__10666),
            .in1(N__16732),
            .in2(N__11053),
            .in3(N__10654),
            .lcout(\uu2.w_addr_displaying_RNI0NG56Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_5_4_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_4_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_5_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13809),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__20942));
    defparam \uu2.trig_rd_det_1_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_5_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10636),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__20942));
    defparam \uu2.trig_rd_det_0_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_5_4_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__14357),
            .in2(_gnd_net_),
            .in3(N__14322),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__20942));
    defparam \buart.Z_rx.hh_0_LC_5_4_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_5_4_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_5_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10624),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__20942));
    defparam \uu0.sec_clkD_LC_5_5_0 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_5_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.sec_clkD_LC_5_5_0  (
            .in0(N__13559),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uu0_sec_clkD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22311),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_5_5_1 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_5_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__11268),
            .in2(_gnd_net_),
            .in3(N__13558),
            .lcout(oneSecStrb),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_5_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_5_5_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_5_5_6  (
            .in0(N__18260),
            .in1(N__18356),
            .in2(N__18455),
            .in3(N__12490),
            .lcout(\Lab_UT.dispString.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_5_5_7 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_5_5_7 .LUT_INIT=16'b0010111110101111;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_5_5_7  (
            .in0(N__11487),
            .in1(N__11464),
            .in2(N__22357),
            .in3(N__11443),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_0_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14260),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22303),
            .ce(N__12316),
            .sr(N__20935));
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_1_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20184),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22303),
            .ce(N__12316),
            .sr(N__20935));
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_2_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20337),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22303),
            .ce(N__12316),
            .sr(N__20935));
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_3_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20522),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22303),
            .ce(N__12316),
            .sr(N__20935));
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_5_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_5_7_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIH15E_2_LC_5_7_1  (
            .in0(N__18426),
            .in1(N__18244),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dispString.un42_dOutP_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_1_LC_5_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_5_7_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_5_7_3  (
            .in0(N__18428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18350),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22294),
            .ce(),
            .sr(N__20933));
    defparam \Lab_UT.dispString.cnt_0_LC_5_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_5_7_4 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_5_7_4  (
            .in0(N__18349),
            .in1(N__11657),
            .in2(N__18261),
            .in3(N__18427),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22294),
            .ce(),
            .sr(N__20933));
    defparam \Lab_UT.didp.ce_0_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_5_7_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_5_7_5  (
            .in0(N__11656),
            .in1(N__17788),
            .in2(_gnd_net_),
            .in3(N__21287),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22294),
            .ce(),
            .sr(N__20933));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_7_6 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_5_7_6  (
            .in0(N__11774),
            .in1(N__12285),
            .in2(N__12604),
            .in3(N__14153),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_7 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__11687),
            .in2(N__10669),
            .in3(N__17396),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_3_LC_5_8_0 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_3_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_3_LC_5_8_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.un1_w_user_cr_3_LC_5_8_0  (
            .in0(N__10754),
            .in1(N__10886),
            .in2(_gnd_net_),
            .in3(N__11702),
            .lcout(\uu2.un1_w_user_crZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_5_8_1  (
            .in0(N__11703),
            .in1(N__10755),
            .in2(N__10698),
            .in3(N__10776),
            .lcout(),
            .ltout(\uu2.un1_w_user_lfZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un20_w_addr_user_1_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.un20_w_addr_user_1_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un20_w_addr_user_1_LC_5_8_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \uu2.un20_w_addr_user_1_LC_5_8_2  (
            .in0(N__10717),
            .in1(N__11459),
            .in2(N__10798),
            .in3(N__11438),
            .lcout(\uu2.un20_w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.un1_w_user_cr_4_LC_5_8_3  (
            .in0(N__11504),
            .in1(N__10685),
            .in2(N__10740),
            .in3(N__10775),
            .lcout(\uu2.un1_w_user_crZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_5_8_4  (
            .in0(N__18358),
            .in1(N__18267),
            .in2(_gnd_net_),
            .in3(N__10858),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22287),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uu2.un1_w_user_lf_3_LC_5_8_5  (
            .in0(N__10887),
            .in1(_gnd_net_),
            .in2(N__11508),
            .in3(N__10733),
            .lcout(\uu2.un1_w_user_lfZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_8_6 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_8_6  (
            .in0(N__18357),
            .in1(_gnd_net_),
            .in2(N__18448),
            .in3(N__18265),
            .lcout(\Lab_UT.dispString.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_8_7 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_5_8_7  (
            .in0(N__18266),
            .in1(N__11776),
            .in2(N__10711),
            .in3(N__13361),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_5_9_0 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_5_9_0  (
            .in0(N__11567),
            .in1(N__18362),
            .in2(N__11254),
            .in3(N__10870),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22279),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_9_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_5_9_1  (
            .in0(N__18361),
            .in1(N__11566),
            .in2(N__11287),
            .in3(N__10914),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_5_9_2 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_5_9_2  (
            .in0(N__10903),
            .in1(N__11747),
            .in2(N__10897),
            .in3(N__13424),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22279),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_3 .LUT_INIT=16'b1100100011111111;
    LogicCell40 \Lab_UT.alarmchar_latch_0_LC_5_9_3  (
            .in0(N__11532),
            .in1(N__11353),
            .in2(N__21041),
            .in3(N__11413),
            .lcout(G_186),
            .ltout(G_186_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_9_4 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_5_9_4  (
            .in0(N__18447),
            .in1(_gnd_net_),
            .in2(N__10873),
            .in3(N__18359),
            .lcout(\Lab_UT.dispString.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_4_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_4_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_4_LC_5_9_5 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \Lab_UT.alarmchar_latch_4_LC_5_9_5  (
            .in0(N__10869),
            .in1(N__10977),
            .in2(N__21042),
            .in3(N__11354),
            .lcout(G_187),
            .ltout(G_187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_6  (
            .in0(N__11565),
            .in1(N__11250),
            .in2(N__10861),
            .in3(N__18360),
            .lcout(\Lab_UT.dispString.dOutP_1_iv_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_5_10_0 .LUT_INIT=16'b0000000001001111;
    LogicCell40 \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_5_10_0  (
            .in0(N__10966),
            .in1(N__10941),
            .in2(N__10981),
            .in3(N__12396),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.justentered_latch_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.justentered_latch_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.justentered_latch_LC_5_10_1 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \Lab_UT.dictrl.justentered_latch_LC_5_10_1  (
            .in0(N__12395),
            .in1(N__10964),
            .in2(N__10852),
            .in3(N__21040),
            .lcout(G_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_10_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_10_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m1_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m1_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m1_LC_5_10_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.m1_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__11352),
            .in2(_gnd_net_),
            .in3(N__11412),
            .lcout(G_182),
            .ltout(G_182_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_5_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_5_10_6 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_5_10_6  (
            .in0(N__10965),
            .in1(N__10940),
            .in2(N__10954),
            .in3(N__12394),
            .lcout(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_7_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_7_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_7_LC_5_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g1_7_LC_5_11_0  (
            .in0(N__15378),
            .in1(N__15558),
            .in2(N__12956),
            .in3(N__12865),
            .lcout(\Lab_UT.dictrl.g1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_5_11_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_3_LC_5_11_1  (
            .in0(N__15698),
            .in1(N__12933),
            .in2(N__20028),
            .in3(N__15377),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_LC_5_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_LC_5_11_2  (
            .in0(N__15553),
            .in1(N__12864),
            .in2(N__10945),
            .in3(N__19578),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_1_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_1_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_1_LC_5_11_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.dictrl.g1_0_1_LC_5_11_3  (
            .in0(N__15699),
            .in1(_gnd_net_),
            .in2(N__20029),
            .in3(N__15554),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_5_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_5_11_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_5_11_4  (
            .in0(N__20127),
            .in1(N__11806),
            .in2(N__10927),
            .in3(N__15194),
            .lcout(\Lab_UT.dictrl.g1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_0_LC_5_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_0_LC_5_11_5 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g2_0_LC_5_11_5  (
            .in0(N__20441),
            .in1(N__20126),
            .in2(_gnd_net_),
            .in3(N__20303),
            .lcout(\Lab_UT.dictrl.g2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_1_LC_5_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_1_LC_5_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_1_LC_5_11_6  (
            .in0(N__12937),
            .in1(N__20442),
            .in2(N__15565),
            .in3(N__12866),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_5_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_5_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_5_11_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_5_11_7  (
            .in0(N__11785),
            .in1(N__10924),
            .in2(N__10918),
            .in3(N__21439),
            .lcout(\Lab_UT.dictrl.N_55_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15563),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__15479),
            .sr(N__20966));
    defparam \buart.Z_rx.shifter_4_LC_5_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12893),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__15479),
            .sr(N__20966));
    defparam \buart.Z_rx.shifter_5_LC_5_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12962),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__15479),
            .sr(N__20966));
    defparam \buart.Z_rx.shifter_3_LC_5_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15389),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__15479),
            .sr(N__20966));
    defparam \buart.Z_rx.shifter_2_rep1_LC_5_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20459),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22268),
            .ce(N__15478),
            .sr(N__20967));
    defparam \buart.Z_rx.shifter_3_rep2_LC_5_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep2_LC_5_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15390),
            .lcout(bu_rx_data_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22268),
            .ce(N__15478),
            .sr(N__20967));
    defparam \buart.Z_rx.shifter_fast_2_LC_5_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_5_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20460),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22268),
            .ce(N__15478),
            .sr(N__20967));
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12963),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22266),
            .ce(N__15476),
            .sr(N__20968));
    defparam \buart.Z_rx.shifter_0_rep1_LC_5_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_rep1_LC_5_14_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__20155),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22266),
            .ce(N__15476),
            .sr(N__20968));
    defparam \buart.Z_rx.shifter_3_rep1_LC_5_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15403),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22266),
            .ce(N__15476),
            .sr(N__20968));
    defparam \buart.Z_rx.shifter_fast_3_LC_5_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_5_15_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__15404),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(N__15475),
            .sr(N__20970));
    defparam \uu2.w_addr_user_2_LC_6_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_6_1_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_2_LC_6_1_0  (
            .in0(N__21945),
            .in1(N__15966),
            .in2(N__20743),
            .in3(N__11000),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_user_1_LC_6_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_6_1_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_user_1_LC_6_1_1  (
            .in0(N__10998),
            .in1(N__15962),
            .in2(_gnd_net_),
            .in3(N__20738),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_user_0_LC_6_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_6_1_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_user_0_LC_6_1_2  (
            .in0(N__15961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10997),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_user_4_LC_6_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_6_1_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_user_4_LC_6_1_3  (
            .in0(N__10999),
            .in1(N__15923),
            .in2(_gnd_net_),
            .in3(N__16185),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_user_5_LC_6_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_6_1_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_5_LC_6_1_4  (
            .in0(N__16186),
            .in1(N__15439),
            .in2(N__15928),
            .in3(N__11001),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_user_6_LC_6_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_6_1_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_6_1_5  (
            .in0(N__11002),
            .in1(N__15927),
            .in2(N__15904),
            .in3(N__16051),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15834));
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6  (
            .in0(_gnd_net_),
            .in1(N__21022),
            .in2(_gnd_net_),
            .in3(N__13932),
            .lcout(\uu2.N_33_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_6_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_6_2_0 .LUT_INIT=16'b0100000110111110;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_6_2_0  (
            .in0(N__13160),
            .in1(N__16251),
            .in2(N__16467),
            .in3(N__11987),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_6_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_6_2_1 .LUT_INIT=16'b0000100101000010;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_6_2_1  (
            .in0(N__11131),
            .in1(N__16119),
            .in2(N__11038),
            .in3(N__11028),
            .lcout(\uu2.bitmap_pmux_sn_i5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_6_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_6_2_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_6_2_2  (
            .in0(N__13159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12097),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_6_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_6_2_3 .LUT_INIT=16'b0001001100010010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_6_2_3  (
            .in0(N__11988),
            .in1(N__16331),
            .in2(N__12106),
            .in3(N__16462),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_N_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_6_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_6_2_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__16429),
            .in2(N__11017),
            .in3(N__11953),
            .lcout(\uu2.N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_6_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_6_2_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_LC_6_2_5  (
            .in0(N__12101),
            .in1(_gnd_net_),
            .in2(N__16262),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__13261),
            .sr(N__20899));
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_6_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_6_2_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_1_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__16255),
            .in2(_gnd_net_),
            .in3(N__12102),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__13261),
            .sr(N__20899));
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_2_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_nesr_1_LC_6_2_7  (
            .in0(N__12103),
            .in1(_gnd_net_),
            .in2(N__16263),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__13261),
            .sr(N__20899));
    defparam \uu2.bitmap_197_LC_6_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_6_3_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_197_LC_6_3_0  (
            .in0(N__17374),
            .in1(N__16564),
            .in2(N__16387),
            .in3(N__16420),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20896));
    defparam \uu2.bitmap_RNITSCU1_69_LC_6_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNITSCU1_69_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNITSCU1_69_LC_6_3_1 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \uu2.bitmap_RNITSCU1_69_LC_6_3_1  (
            .in0(N__11008),
            .in1(N__16345),
            .in2(N__11129),
            .in3(N__16513),
            .lcout(\uu2.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_6_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_6_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_0_LC_6_3_2  (
            .in0(N__13953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11110),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20896));
    defparam \uu2.w_addr_displaying_fast_2_LC_6_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_6_3_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_6_3_3  (
            .in0(N__11112),
            .in1(N__13957),
            .in2(N__20703),
            .in3(N__11989),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20896));
    defparam \uu2.w_addr_displaying_2_LC_6_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_6_3_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_2_LC_6_3_4  (
            .in0(N__20681),
            .in1(N__11111),
            .in2(N__13960),
            .in3(N__21776),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20896));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_3_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_3_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_3_5  (
            .in0(N__21775),
            .in1(N__16112),
            .in2(N__11130),
            .in3(N__20680),
            .lcout(\uu2.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_6_3_6 .LUT_INIT=16'b1000000100000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_6_3_6  (
            .in0(N__16111),
            .in1(N__21774),
            .in2(N__11128),
            .in3(N__11848),
            .lcout(\uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_3_7 .LUT_INIT=16'b0110101000001000;
    LogicCell40 \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_3_7  (
            .in0(N__21773),
            .in1(N__20679),
            .in2(N__16128),
            .in3(N__13175),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_3_LC_6_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_6_4_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_6_4_0  (
            .in0(N__12122),
            .in1(N__17142),
            .in2(_gnd_net_),
            .in3(N__11192),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(),
            .sr(N__20945));
    defparam \Lab_UT.didp.ce_1_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_6_4_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_6_4_1  (
            .in0(N__13469),
            .in1(N__11169),
            .in2(N__11654),
            .in3(N__17604),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(),
            .sr(N__20945));
    defparam \Lab_UT.didp.reset_0_LC_6_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_6_4_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_6_4_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_6_4_2  (
            .in0(N__17605),
            .in1(N__13470),
            .in2(N__11173),
            .in3(N__11637),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(),
            .sr(N__20945));
    defparam \Lab_UT.didp.reset_2_LC_6_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_6_4_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_6_4_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_6_4_4  (
            .in0(N__12123),
            .in1(N__17143),
            .in2(_gnd_net_),
            .in3(N__11193),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(),
            .sr(N__20945));
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_4_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_4_5  (
            .in0(N__13468),
            .in1(N__11168),
            .in2(N__11653),
            .in3(N__17603),
            .lcout(\Lab_UT.didp.ce_12_1 ),
            .ltout(\Lab_UT.didp.ce_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_4_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_4_6  (
            .in0(N__12121),
            .in1(_gnd_net_),
            .in2(N__11179),
            .in3(N__17141),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_6_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_6_4_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_6_4_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_6_4_7  (
            .in0(N__13849),
            .in1(N__17440),
            .in2(N__11176),
            .in3(N__17050),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(),
            .sr(N__20945));
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_6_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_6_5_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNIBN0Q1_2_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__11229),
            .in2(_gnd_net_),
            .in3(N__16956),
            .lcout(\Lab_UT.didp.un1_dicLdMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_6_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_6_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__17717),
            .in2(_gnd_net_),
            .in3(N__17277),
            .lcout(\Lab_UT.didp.countrce1.ce_12_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_5_2  (
            .in0(N__17278),
            .in1(N__17721),
            .in2(_gnd_net_),
            .in3(N__17602),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_5_3 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_5_3  (
            .in0(N__17646),
            .in1(N__13462),
            .in2(N__11158),
            .in3(N__20511),
            .lcout(\Lab_UT.didp.countrce1.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_6_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_2_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__16994),
            .in2(_gnd_net_),
            .in3(N__17941),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_6_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_6_5_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_6_5_5  (
            .in0(N__16955),
            .in1(N__20336),
            .in2(N__11155),
            .in3(N__17225),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_6_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_6_5_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_6_5_6  (
            .in0(N__17226),
            .in1(N__17992),
            .in2(N__11152),
            .in3(N__17952),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22298),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_5_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_5_7  (
            .in0(N__16995),
            .in1(N__16954),
            .in2(_gnd_net_),
            .in3(N__14265),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_6_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_6_6_0  (
            .in0(N__13463),
            .in1(N__17302),
            .in2(N__17764),
            .in3(N__11296),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22290),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_6_1 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_6_1  (
            .in0(N__13425),
            .in1(N__17045),
            .in2(N__13464),
            .in3(N__13826),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_6_2 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_3_LC_6_6_2  (
            .in0(N__13827),
            .in1(N__11686),
            .in2(N__11655),
            .in3(N__18433),
            .lcout(\Lab_UT.dispString.N_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_6_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__18248),
            .in2(_gnd_net_),
            .in3(N__18319),
            .lcout(\Lab_UT.dispString.N_143 ),
            .ltout(\Lab_UT.dispString.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_6_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_6_6_4 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIKUO21_1_LC_6_6_4  (
            .in0(N__11272),
            .in1(N__13564),
            .in2(N__11257),
            .in3(N__18432),
            .lcout(\Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_6_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_6_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dispString.rdy_LC_6_6_5  (
            .in0(N__18434),
            .in1(N__11641),
            .in2(N__18268),
            .in3(N__18320),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22290),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_6_7 .LUT_INIT=16'b0000111000000001;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_6_6_7  (
            .in0(N__16957),
            .in1(N__11233),
            .in2(N__18013),
            .in3(N__11212),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22290),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_6_7_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_6_7_0  (
            .in0(N__16996),
            .in1(N__14438),
            .in2(N__12226),
            .in3(N__13871),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_6_7_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_6_7_1  (
            .in0(N__18415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18242),
            .lcout(\Lab_UT.dispString.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_6_7_2 .LUT_INIT=16'b0010001001000101;
    LogicCell40 \Lab_UT.dispString.cnt_RNIKUO21_2_LC_6_7_2  (
            .in0(N__18243),
            .in1(N__18417),
            .in2(N__11665),
            .in3(N__18325),
            .lcout(\Lab_UT.dispString.N_102 ),
            .ltout(\Lab_UT.dispString.N_102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_7_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_6_7_3  (
            .in0(N__18326),
            .in1(N__11573),
            .in2(N__11539),
            .in3(N__11536),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_6_7_4 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_6_7_4  (
            .in0(N__11748),
            .in1(N__11521),
            .in2(N__11515),
            .in3(N__14400),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22283),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_7_5 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_7_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \uu2.un4_w_user_data_rdy_0_LC_6_7_5  (
            .in0(N__11477),
            .in1(N__11460),
            .in2(_gnd_net_),
            .in3(N__11439),
            .lcout(\uu2.un4_w_user_data_rdyZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_6_7_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIFV4E_1_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__18416),
            .in2(_gnd_net_),
            .in3(N__18324),
            .lcout(\Lab_UT.dispString.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_6_7_7 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \Lab_UT.didp.ce_RNIHGGI1_3_LC_6_7_7  (
            .in0(N__17121),
            .in1(_gnd_net_),
            .in2(N__12339),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.un1_dicLdMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_8_0 .LUT_INIT=16'b0000100000000010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_8_0  (
            .in0(N__11422),
            .in1(N__17188),
            .in2(N__11365),
            .in3(N__13372),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_1 .LUT_INIT=16'b1000000001000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_1  (
            .in0(N__17728),
            .in1(N__11305),
            .in2(N__11299),
            .in3(N__13392),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_8_3 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_6_8_3  (
            .in0(N__11775),
            .in1(N__12225),
            .in2(N__13879),
            .in3(N__11688),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_8_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_6_8_4  (
            .in0(N__12603),
            .in1(N__11758),
            .in2(N__11752),
            .in3(N__12368),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_6_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_6_8_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_6_8_5  (
            .in0(N__11749),
            .in1(N__11722),
            .in2(N__11716),
            .in3(N__13391),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_8_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_6_8_6  (
            .in0(N__11689),
            .in1(N__12580),
            .in2(N__11664),
            .in3(N__16590),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_0_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14253),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22272),
            .ce(N__11587),
            .sr(N__20936));
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_1_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20169),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22272),
            .ce(N__11587),
            .sr(N__20936));
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_2_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20325),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22272),
            .ce(N__11587),
            .sr(N__20936));
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_3_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20487),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22272),
            .ce(N__11587),
            .sr(N__20936));
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_0_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14257),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22270),
            .ce(N__12574),
            .sr(N__20938));
    defparam \Lab_UT.dictrl.g1_8_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_8_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_8_LC_6_11_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.g1_8_LC_6_11_0  (
            .in0(N__19457),
            .in1(N__19735),
            .in2(N__15785),
            .in3(N__15708),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_6_11_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_6_11_1  (
            .in0(N__21438),
            .in1(N__11800),
            .in2(N__11791),
            .in3(N__19905),
            .lcout(\Lab_UT.dictrl.G_14_0_a2_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_11_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_11_2  (
            .in0(N__19906),
            .in1(N__21437),
            .in2(_gnd_net_),
            .in3(N__12952),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_25_i_o3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_11_3 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_11_3  (
            .in0(N__20312),
            .in1(N__20452),
            .in2(N__11788),
            .in3(N__20177),
            .lcout(\Lab_UT.dictrl.G_25_i_o3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_11_5 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_11_5  (
            .in0(N__20311),
            .in1(N__20631),
            .in2(N__20162),
            .in3(N__15388),
            .lcout(\Lab_UT.dictrl.g0_5_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_11_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.g0_6_1_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__12883),
            .in2(_gnd_net_),
            .in3(N__12951),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_11_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_11_7  (
            .in0(N__20632),
            .in1(N__15564),
            .in2(N__11779),
            .in3(N__15387),
            .lcout(\Lab_UT.dictrl.g0_6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_12_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m37_N_2L1_LC_6_12_0  (
            .in0(N__14219),
            .in1(N__12867),
            .in2(N__20301),
            .in3(N__19991),
            .lcout(\Lab_UT.dictrl.m37_N_2LZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__20261),
            .in2(_gnd_net_),
            .in3(N__14220),
            .lcout(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_6_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_1_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__12990),
            .in2(_gnd_net_),
            .in3(N__13022),
            .lcout(\Lab_UT.dictrl.m13_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_4_LC_6_12_3 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_6_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \resetGen.escKey_4_LC_6_12_3  (
            .in0(N__15386),
            .in1(N__20183),
            .in2(N__20483),
            .in3(N__14221),
            .lcout(),
            .ltout(\resetGen.escKeyZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_6_12_4 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_6_12_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \resetGen.escKey_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__11812),
            .in2(N__11839),
            .in3(N__18078),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_5_LC_6_12_5 .C_ON=1'b0;
    defparam \resetGen.escKey_5_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_5_LC_6_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \resetGen.escKey_5_LC_6_12_5  (
            .in0(N__15561),
            .in1(N__12950),
            .in2(N__12885),
            .in3(N__20262),
            .lcout(\resetGen.escKeyZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_12_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_5_LC_6_12_6  (
            .in0(N__12949),
            .in1(N__12868),
            .in2(N__15787),
            .in3(N__15384),
            .lcout(\Lab_UT.dictrl.g1_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_6_12_7 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_5_LC_6_12_7  (
            .in0(N__15385),
            .in1(N__15562),
            .in2(N__21289),
            .in3(N__12884),
            .lcout(\Lab_UT.dictrl.G_25_i_o3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_6_13_0 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_6_13_0  (
            .in0(N__19990),
            .in1(N__13028),
            .in2(N__19920),
            .in3(N__12992),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_1_LC_6_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_6_13_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_6_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20274),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22265),
            .ce(N__15477),
            .sr(N__20969));
    defparam \buart.Z_rx.shifter_1_rep1_LC_6_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_6_13_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_6_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_6_13_2  (
            .in0(N__20275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22265),
            .ce(N__15477),
            .sr(N__20969));
    defparam \buart.Z_rx.shifter_2_LC_6_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_6_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_6_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20461),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22265),
            .ce(N__15477),
            .sr(N__20969));
    defparam \Lab_UT.dictrl.g1_1_5_LC_6_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_5_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_5_LC_6_14_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.g1_1_5_LC_6_14_2  (
            .in0(N__13024),
            .in1(N__11910),
            .in2(N__15327),
            .in3(N__15646),
            .lcout(\Lab_UT.dictrl.g1_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_6_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_6_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_6_14_5  (
            .in0(N__12825),
            .in1(N__14689),
            .in2(N__11911),
            .in3(N__13023),
            .lcout(\Lab_UT.dictrl.g1_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m34_1_LC_6_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m34_1_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m34_1_LC_6_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m34_1_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__12991),
            .in2(_gnd_net_),
            .in3(N__15645),
            .lcout(\Lab_UT.dictrl.m34Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_8_LC_7_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_8_LC_7_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_8_LC_7_1_0 .LUT_INIT=16'b1111101100000100;
    LogicCell40 \uu2.w_addr_displaying_fast_8_LC_7_1_0  (
            .in0(N__12796),
            .in1(N__13947),
            .in2(N__11895),
            .in3(N__16759),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20902));
    defparam \uu2.w_addr_displaying_8_LC_7_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_7_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_7_1_1 .LUT_INIT=16'b1100110011000110;
    LogicCell40 \uu2.w_addr_displaying_8_LC_7_1_1  (
            .in0(N__13945),
            .in1(N__13312),
            .in2(N__12811),
            .in3(N__11886),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20902));
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_7_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_7_1_2 .LUT_INIT=16'b0000001011111111;
    LogicCell40 \uu2.w_addr_displaying_RNI0ES07_8_LC_7_1_2  (
            .in0(N__13311),
            .in1(N__12804),
            .in2(N__11893),
            .in3(N__21866),
            .lcout(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ),
            .ltout(\uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_7_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_7_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_7_1_3 .LUT_INIT=16'b1100111100110000;
    LogicCell40 \uu2.w_addr_displaying_4_LC_7_1_3  (
            .in0(_gnd_net_),
            .in1(N__11882),
            .in2(N__11899),
            .in3(N__13173),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20902));
    defparam \uu2.w_addr_displaying_5_LC_7_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_7_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_7_1_4 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_7_1_4  (
            .in0(N__13174),
            .in1(N__13946),
            .in2(N__11894),
            .in3(N__13102),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20902));
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_7_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_7_1_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNO_0_6_LC_7_1_5  (
            .in0(N__13101),
            .in1(N__11881),
            .in2(_gnd_net_),
            .in3(N__13172),
            .lcout(\uu2.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_7_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_7_1_6 .LUT_INIT=16'b0001010000011000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_7_1_6  (
            .in0(N__13214),
            .in1(N__16311),
            .in2(N__13326),
            .in3(N__13099),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_7_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_7_1_7 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_7_1_7  (
            .in0(N__13100),
            .in1(N__13310),
            .in2(N__16325),
            .in3(N__13215),
            .lcout(\uu2.bitmap_pmux_sn_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_7_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_7_2_1 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_40_LC_7_2_1  (
            .in0(N__14667),
            .in1(N__14502),
            .in2(N__14628),
            .in3(N__14576),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__20901));
    defparam \uu2.bitmap_75_LC_7_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_7_2_2 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_75_LC_7_2_2  (
            .in0(N__14577),
            .in1(N__14621),
            .in2(N__14506),
            .in3(N__14668),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__20901));
    defparam \uu2.bitmap_203_LC_7_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_7_2_3 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_203_LC_7_2_3  (
            .in0(N__14666),
            .in1(N__14501),
            .in2(N__14627),
            .in3(N__14575),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__20901));
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_4 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_4  (
            .in0(N__11986),
            .in1(N__11945),
            .in2(_gnd_net_),
            .in3(N__11968),
            .lcout(\uu2.bitmap_pmux_sn_N_54_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.bitmap_RNIJS4P_162_LC_7_2_5  (
            .in0(N__11946),
            .in1(N__16501),
            .in2(_gnd_net_),
            .in3(N__13477),
            .lcout(),
            .ltout(\uu2.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6  (
            .in0(_gnd_net_),
            .in1(N__13522),
            .in2(N__11962),
            .in3(N__11959),
            .lcout(\uu2.bitmap_RNI2Q8F1Z0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \uu2.bitmap_RNIBPBO_40_LC_7_2_7  (
            .in0(N__11944),
            .in1(N__11917),
            .in2(N__13486),
            .in3(N__16761),
            .lcout(\uu2.bitmap_pmux_26_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_7_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_7_3_0 .LUT_INIT=16'b0110011100011111;
    LogicCell40 \uu2.bitmap_93_LC_7_3_0  (
            .in0(N__16835),
            .in1(N__16881),
            .in2(N__16810),
            .in3(N__16912),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__20900));
    defparam \uu2.bitmap_221_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_7_3_1 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \uu2.bitmap_221_LC_7_3_1  (
            .in0(N__16911),
            .in1(N__16806),
            .in2(N__16885),
            .in3(N__16834),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__20900));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_7_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_7_3_2  (
            .in0(N__16234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12105),
            .lcout(\uu2.N_31_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI6MCU1_93_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI6MCU1_93_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI6MCU1_93_LC_7_3_3 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \uu2.bitmap_RNI6MCU1_93_LC_7_3_3  (
            .in0(N__12073),
            .in1(N__16236),
            .in2(N__12067),
            .in3(N__16198),
            .lcout(\uu2.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIPIHG1_75_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_7_3_4 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.bitmap_RNIPIHG1_75_LC_7_3_4  (
            .in0(N__16235),
            .in1(N__12055),
            .in2(N__12049),
            .in3(N__13969),
            .lcout(),
            .ltout(\uu2.N_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_7_3_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_7_3_5  (
            .in0(N__16138),
            .in1(N__12036),
            .in2(N__12040),
            .in3(N__12139),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_27_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI72CH8_69_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI72CH8_69_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI72CH8_69_LC_7_3_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.bitmap_RNI72CH8_69_LC_7_3_6  (
            .in0(N__12037),
            .in1(N__12028),
            .in2(N__12022),
            .in3(N__12019),
            .lcout(\uu2.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_7_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_7_4_0 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_308_LC_7_4_0  (
            .in0(N__14025),
            .in1(N__14062),
            .in2(N__14131),
            .in3(N__14091),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_212_LC_7_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_7_4_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_212_LC_7_4_1  (
            .in0(N__14090),
            .in1(N__14117),
            .in2(N__14068),
            .in3(N__14024),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_84_LC_7_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_7_4_2 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_84_LC_7_4_2  (
            .in0(N__14027),
            .in1(N__14064),
            .in2(N__14133),
            .in3(N__14093),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_180_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_7_4_3 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_180_LC_7_4_3  (
            .in0(N__14089),
            .in1(N__14116),
            .in2(N__14067),
            .in3(N__14023),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_52_LC_7_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_7_4_4 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_52_LC_7_4_4  (
            .in0(N__14026),
            .in1(N__14063),
            .in2(N__14132),
            .in3(N__14092),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIB3QK_52_LC_7_4_5  (
            .in0(N__16760),
            .in1(N__12178),
            .in2(_gnd_net_),
            .in3(N__12172),
            .lcout(\uu2.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_7_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_7_4_6 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_87_LC_7_4_6  (
            .in0(N__14028),
            .in1(N__14065),
            .in2(N__14134),
            .in3(N__14094),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20897));
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \uu2.bitmap_RNIRMQA1_84_LC_7_4_7  (
            .in0(N__12154),
            .in1(N__13990),
            .in2(N__12148),
            .in3(N__16717),
            .lcout(\uu2.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_5_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_5_0  (
            .in0(N__13602),
            .in1(N__14297),
            .in2(N__12256),
            .in3(N__12457),
            .lcout(\Lab_UT.didp.un24_ce_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_5_1 .LUT_INIT=16'b0000001000001101;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_7_5_1  (
            .in0(N__17889),
            .in1(N__16671),
            .in2(N__12523),
            .in3(N__14164),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22312),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_2  (
            .in0(N__17520),
            .in1(N__14296),
            .in2(_gnd_net_),
            .in3(N__12373),
            .lcout(\Lab_UT.sec1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_5_3 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_5_3  (
            .in0(N__13570),
            .in1(N__20339),
            .in2(N__17895),
            .in3(N__12253),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_5_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_7_5_4  (
            .in0(N__12254),
            .in1(N__12519),
            .in2(N__12301),
            .in3(N__16650),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22312),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_7_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_7_5_5  (
            .in0(N__12286),
            .in1(N__12248),
            .in2(_gnd_net_),
            .in3(N__17521),
            .lcout(\Lab_UT.sec1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_6  (
            .in0(N__17519),
            .in1(N__12456),
            .in2(_gnd_net_),
            .in3(N__12489),
            .lcout(\Lab_UT.sec1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_5_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_5_7  (
            .in0(N__14298),
            .in1(N__12252),
            .in2(_gnd_net_),
            .in3(N__13601),
            .lcout(\Lab_UT.didp.countrce2.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_1 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_1  (
            .in0(N__12298),
            .in1(N__20523),
            .in2(N__17896),
            .in3(N__12458),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_7_6_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_7_6_2  (
            .in0(N__16657),
            .in1(N__12459),
            .in2(N__12289),
            .in3(N__12517),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22304),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_6_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_6_3  (
            .in0(N__17578),
            .in1(N__12281),
            .in2(N__12255),
            .in3(N__13631),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_7_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_7_6_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_7_6_4  (
            .in0(N__17397),
            .in1(N__14532),
            .in2(N__17940),
            .in3(N__17429),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_6_5  (
            .in0(N__16985),
            .in1(N__12224),
            .in2(_gnd_net_),
            .in3(N__17510),
            .lcout(\Lab_UT.min2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_6 .LUT_INIT=16'b1100001101010101;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_6  (
            .in0(N__20187),
            .in1(N__14301),
            .in2(N__13609),
            .in3(N__17894),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_6_7 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_7_6_7  (
            .in0(N__12518),
            .in1(N__13606),
            .in2(N__12493),
            .in3(N__16656),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22304),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_7_7_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_7_7_0  (
            .in0(N__13662),
            .in1(N__12482),
            .in2(N__12460),
            .in3(N__13595),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_7_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_7_7_1  (
            .in0(N__14374),
            .in1(N__12430),
            .in2(N__12424),
            .in3(N__12421),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_7_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_7_7_2  (
            .in0(N__12349),
            .in1(N__12415),
            .in2(N__12406),
            .in3(N__12403),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_7_7_3 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_7_7_3  (
            .in0(N__12369),
            .in1(N__17227),
            .in2(N__14305),
            .in3(N__14154),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_7_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_7_4  (
            .in0(N__17109),
            .in1(N__14437),
            .in2(_gnd_net_),
            .in3(N__14264),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_7_5 .LUT_INIT=16'b0101000001000001;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_7_7_5  (
            .in0(N__14746),
            .in1(N__17110),
            .in2(N__12343),
            .in3(N__12340),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_0  (
            .in0(N__21251),
            .in1(N__20615),
            .in2(N__18949),
            .in3(N__21025),
            .lcout(\Lab_UT.didp.regrce4.LdAMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_7_8_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_1_LC_7_8_1  (
            .in0(N__18368),
            .in1(N__18252),
            .in2(N__18456),
            .in3(N__14531),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_8_2 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_7_8_2  (
            .in0(N__12599),
            .in1(N__18369),
            .in2(N__12583),
            .in3(N__13661),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_8_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__14809),
            .in2(_gnd_net_),
            .in3(N__21024),
            .lcout(\Lab_UT.didp.regrce1.LdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20170),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__12567),
            .sr(N__20939));
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20330),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__12567),
            .sr(N__20939));
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20515),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__12567),
            .sr(N__20939));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_10_0 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_10_0  (
            .in0(N__19053),
            .in1(N__15223),
            .in2(N__15198),
            .in3(N__13048),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_10_1 .LUT_INIT=16'b1110111000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_10_1  (
            .in0(N__12547),
            .in1(N__12535),
            .in2(N__12529),
            .in3(N__21166),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_10_2 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_10_2  (
            .in0(N__19258),
            .in1(N__18066),
            .in2(N__12526),
            .in3(N__12637),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_25_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_3 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_LC_7_10_3  (
            .in0(N__18157),
            .in1(N__17824),
            .in2(N__12640),
            .in3(N__12631),
            .lcout(\Lab_UT.un1_next_state66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22275),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_4 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_4  (
            .in0(N__19256),
            .in1(N__18065),
            .in2(N__18741),
            .in3(N__12724),
            .lcout(\Lab_UT.dictrl.G_25_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6  (
            .in0(N__21167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19052),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_7 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_7  (
            .in0(N__18067),
            .in1(N__19257),
            .in2(N__18601),
            .in3(N__21058),
            .lcout(\Lab_UT.dictrl.G_25_i_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_11_0 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_11_0  (
            .in0(N__19822),
            .in1(N__20037),
            .in2(N__19919),
            .in3(N__19588),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_18_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_11_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_11_1  (
            .in0(N__15187),
            .in1(N__12646),
            .in2(N__12625),
            .in3(N__21429),
            .lcout(\Lab_UT.dictrl.N_22_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_11_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_11_2  (
            .in0(N__21428),
            .in1(N__15186),
            .in2(N__18770),
            .in3(N__19636),
            .lcout(\Lab_UT.dictrl.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_11_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_11_3  (
            .in0(N__12673),
            .in1(N__12622),
            .in2(N__12616),
            .in3(N__21430),
            .lcout(\Lab_UT.dictrl.N_57_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_7_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_7_11_4 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_7_11_4  (
            .in0(N__19455),
            .in1(N__19731),
            .in2(_gnd_net_),
            .in3(N__15788),
            .lcout(shifter_1_rep1_RNI0FPF),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_7_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_7_11_5 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_7_11_5  (
            .in0(N__15789),
            .in1(N__19821),
            .in2(N__19738),
            .in3(N__19456),
            .lcout(N_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_7_11_6 .LUT_INIT=16'b0000101001100110;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_7_11_6  (
            .in0(N__21427),
            .in1(N__12661),
            .in2(N__18769),
            .in3(N__21159),
            .lcout(\Lab_UT.dictrl.m19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_2_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_2_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_2_LC_7_11_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.didp.g0_0_2_LC_7_11_7  (
            .in0(N__18046),
            .in1(N__12772),
            .in2(N__19245),
            .in3(N__12715),
            .lcout(\Lab_UT.didp.g0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_0  (
            .in0(N__14223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19908),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_12_1  (
            .in0(N__15259),
            .in1(N__20469),
            .in2(N__12676),
            .in3(N__12740),
            .lcout(\Lab_UT.dictrl.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_7_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_7_12_2  (
            .in0(N__19819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12667),
            .lcout(\Lab_UT.dictrl.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_7_12_3 .LUT_INIT=16'b0000101000101010;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_7_12_3  (
            .in0(N__19907),
            .in1(N__13039),
            .in2(N__19723),
            .in3(N__12994),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_7_12_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_7_12_4  (
            .in0(N__19820),
            .in1(_gnd_net_),
            .in2(N__12655),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m37_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m37_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m37_LC_7_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m37_LC_7_12_5  (
            .in0(N__15559),
            .in1(N__12652),
            .in2(N__15307),
            .in3(N__12957),
            .lcout(\Lab_UT.dictrl.next_state6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_8_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_8_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_8_LC_7_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_8_LC_7_12_6  (
            .in0(N__14222),
            .in1(N__15258),
            .in2(N__12742),
            .in3(N__20033),
            .lcout(\Lab_UT.dictrl.N_72_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m34_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m34_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m34_LC_7_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m34_LC_7_12_7  (
            .in0(N__15560),
            .in1(N__12886),
            .in2(N__15306),
            .in3(N__12958),
            .lcout(\Lab_UT.dictrl.N_67_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_13_0 .LUT_INIT=16'b0011111110101010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_13_0  (
            .in0(N__12748),
            .in1(N__12741),
            .in2(N__15257),
            .in3(N__12763),
            .lcout(),
            .ltout(\Lab_UT.i8_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_13_1 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \Lab_UT.didp.g0_0_2_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__12754),
            .in2(N__12775),
            .in3(N__21168),
            .lcout(\Lab_UT.didp.g0_0_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_13_2  (
            .in0(N__15225),
            .in1(N__20014),
            .in2(N__15715),
            .in3(N__15184),
            .lcout(\Lab_UT.dictrl.g0_0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_13_3  (
            .in0(N__19895),
            .in1(N__21278),
            .in2(_gnd_net_),
            .in3(N__21419),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_13_4 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_13_4  (
            .in0(N__19800),
            .in1(N__20015),
            .in2(N__12757),
            .in3(N__19587),
            .lcout(\Lab_UT.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_13_5  (
            .in0(N__15183),
            .in1(N__19070),
            .in2(_gnd_net_),
            .in3(N__15224),
            .lcout(\Lab_UT.dictrl.g0_0_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_13_6  (
            .in0(N__21169),
            .in1(N__15185),
            .in2(N__21440),
            .in3(N__21288),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.m22_1_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__15783),
            .in2(_gnd_net_),
            .in3(N__19451),
            .lcout(\Lab_UT.dictrl.m22Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_LC_7_14_0 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g2_LC_7_14_0  (
            .in0(N__19695),
            .in1(N__15786),
            .in2(_gnd_net_),
            .in3(N__19452),
            .lcout(\Lab_UT.dictrl.gZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m5_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m5_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m5_LC_7_14_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.m5_LC_7_14_1  (
            .in0(N__12826),
            .in1(N__19365),
            .in2(N__19494),
            .in3(N__15649),
            .lcout(N_63_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_7_14_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_11_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__15624),
            .in2(_gnd_net_),
            .in3(N__19403),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_7_14_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_10_LC_7_14_4  (
            .in0(N__15076),
            .in1(N__19453),
            .in2(N__13051),
            .in3(N__12894),
            .lcout(\Lab_UT.dictrl.N_72_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m7_a0_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m7_a0_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m7_a0_LC_7_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.m7_a0_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__13038),
            .in2(_gnd_net_),
            .in3(N__12993),
            .lcout(m7_a0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_rep1_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12964),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__15473),
            .sr(N__20972));
    defparam \buart.Z_rx.shifter_fast_4_LC_7_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_7_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_7_15_2  (
            .in0(N__12895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__15473),
            .sr(N__20972));
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_7_15_4  (
            .in0(N__15524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__15473),
            .sr(N__20972));
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15599),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__15473),
            .sr(N__20972));
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_8_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_8_1_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_8_1_0  (
            .in0(N__16321),
            .in1(N__13103),
            .in2(N__13224),
            .in3(N__13170),
            .lcout(\uu2.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_6_LC_8_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_8_1_1 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_8_1_1 .LUT_INIT=16'b1111100000001111;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_8_1_1  (
            .in0(N__13325),
            .in1(N__16323),
            .in2(N__13270),
            .in3(N__13220),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_ness_6C_net ),
            .ce(N__13260),
            .sr(N__20905));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_1_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_8_1_2  (
            .in0(N__13219),
            .in1(N__16047),
            .in2(_gnd_net_),
            .in3(N__21901),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_1_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_8_1_3  (
            .in0(N__13171),
            .in1(N__16187),
            .in2(_gnd_net_),
            .in3(N__21899),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_8_1_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_8_1_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_8_1_4  (
            .in0(N__21900),
            .in1(N__15443),
            .in2(_gnd_net_),
            .in3(N__13104),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_8_1_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_8_1_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_8_1_5  (
            .in0(N__15444),
            .in1(N__16188),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.un426_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_8_1_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_8_1_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_8_1_6  (
            .in0(N__16322),
            .in1(N__16013),
            .in2(_gnd_net_),
            .in3(N__21902),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_8_1_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_8_1_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_8_1_7  (
            .in0(N__16014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16050),
            .lcout(\uu2.vbuf_w_addr_user.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_LC_8_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_8_2_0 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uu2.w_addr_displaying_7_LC_8_2_0  (
            .in0(N__13943),
            .in1(N__13896),
            .in2(_gnd_net_),
            .in3(N__16324),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__13944),
            .in2(_gnd_net_),
            .in3(N__16249),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.bitmap_111_LC_8_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_8_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13563),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.vram_rd_clk_det_0_LC_8_2_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_8_2_3 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_8_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14362),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.vram_rd_clk_det_1_LC_8_2_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_8_2_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_8_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13512),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.bitmap_296_LC_8_2_5 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_8_2_5 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_296_LC_8_2_5  (
            .in0(N__14584),
            .in1(N__14609),
            .in2(N__14500),
            .in3(N__14658),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \uu2.bitmap_168_LC_8_2_6 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_8_2_6 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_168_LC_8_2_6  (
            .in0(N__14657),
            .in1(N__14488),
            .in2(N__14622),
            .in3(N__14583),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20903));
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .LUT_INIT=16'b0100010011000000;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_8_3_0  (
            .in0(N__18661),
            .in1(N__21282),
            .in2(N__18634),
            .in3(N__21165),
            .lcout(\Lab_UT.dictrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22333),
            .ce(N__19342),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1  (
            .in0(N__17509),
            .in1(N__13471),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\Lab_UT.sec2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2  (
            .in0(N__17725),
            .in1(N__13393),
            .in2(_gnd_net_),
            .in3(N__17508),
            .lcout(\Lab_UT.sec2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3  (
            .in0(N__17505),
            .in1(_gnd_net_),
            .in2(N__17180),
            .in3(N__13371),
            .lcout(\Lab_UT.min2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4  (
            .in0(N__14451),
            .in1(N__13878),
            .in2(_gnd_net_),
            .in3(N__17507),
            .lcout(\Lab_UT.min1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_3_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_3_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__14452),
            .in2(_gnd_net_),
            .in3(N__16636),
            .lcout(\Lab_UT.didp.reset_12_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6  (
            .in0(N__13837),
            .in1(N__17046),
            .in2(_gnd_net_),
            .in3(N__17506),
            .lcout(\Lab_UT.min1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_8_3_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_8_3_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_8_3_7  (
            .in0(N__13813),
            .in1(N__15585),
            .in2(_gnd_net_),
            .in3(N__13795),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_4_0  (
            .in0(N__13669),
            .in1(N__13607),
            .in2(_gnd_net_),
            .in3(N__17503),
            .lcout(\Lab_UT.sec1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_8_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_8_4_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_8_4_1  (
            .in0(N__17502),
            .in1(N__17591),
            .in2(_gnd_net_),
            .in3(N__13639),
            .lcout(\Lab_UT.sec2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__16635),
            .in2(_gnd_net_),
            .in3(N__14450),
            .lcout(\Lab_UT.didp.countrce4.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_3  (
            .in0(N__13608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14299),
            .lcout(\Lab_UT.didp.countrce2.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_8_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_8_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_8_4_4  (
            .in0(N__14401),
            .in1(N__17271),
            .in2(_gnd_net_),
            .in3(N__17504),
            .lcout(\Lab_UT.sec2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_8_4_5 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \uu2.r_data_rdy_LC_8_4_5  (
            .in0(N__14358),
            .in1(N__14326),
            .in2(N__21043),
            .in3(N__21657),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_4_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_4_6  (
            .in0(N__14300),
            .in1(N__17890),
            .in2(_gnd_net_),
            .in3(N__14266),
            .lcout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_8_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_8_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_8_4_7  (
            .in0(N__17501),
            .in1(N__17235),
            .in2(_gnd_net_),
            .in3(N__14158),
            .lcout(\Lab_UT.min2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_8_5_0 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_8_5_0 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_215_LC_8_5_0  (
            .in0(N__14130),
            .in1(N__14095),
            .in2(N__14066),
            .in3(N__14029),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20898));
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_5_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_5_1 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \uu2.bitmap_RNIOPSS_212_LC_8_5_1  (
            .in0(N__14002),
            .in1(N__13996),
            .in2(N__13984),
            .in3(N__16714),
            .lcout(\uu2.bitmap_pmux_17_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_0_LC_8_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__13958),
            .in2(_gnd_net_),
            .in3(N__13983),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20898));
    defparam \uu2.bitmap_RNI65TM_72_LC_8_5_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI65TM_72_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI65TM_72_LC_8_5_3 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \uu2.bitmap_RNI65TM_72_LC_8_5_3  (
            .in0(N__13982),
            .in1(N__14674),
            .in2(N__14545),
            .in3(N__16715),
            .lcout(\uu2.bitmap_pmux_16_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_7_LC_8_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_5_4 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_8_5_4  (
            .in0(N__16716),
            .in1(N__13959),
            .in2(_gnd_net_),
            .in3(N__13900),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20898));
    defparam \uu2.bitmap_72_LC_8_5_5 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_8_5_5 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_72_LC_8_5_5  (
            .in0(N__14564),
            .in1(N__14626),
            .in2(N__14499),
            .in3(N__14648),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20898));
    defparam \uu2.bitmap_200_LC_8_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_8_5_6 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_200_LC_8_5_6  (
            .in0(N__14647),
            .in1(N__14484),
            .in2(N__14629),
            .in3(N__14563),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20898));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_0  (
            .in0(N__17929),
            .in1(N__17500),
            .in2(_gnd_net_),
            .in3(N__14536),
            .lcout(\Lab_UT.min2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_6_1 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_6_1  (
            .in0(N__16632),
            .in1(N__14433),
            .in2(N__17125),
            .in3(N__20199),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_6_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_8_6_2  (
            .in0(N__14747),
            .in1(N__14773),
            .in2(N__14455),
            .in3(N__16633),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_8_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_8_6_3  (
            .in0(N__16631),
            .in1(N__14432),
            .in2(_gnd_net_),
            .in3(N__17431),
            .lcout(\Lab_UT.didp.countrce4.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_6_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_8_6_4  (
            .in0(N__17044),
            .in1(N__17008),
            .in2(N__14754),
            .in3(N__14772),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_6_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_8_6_5  (
            .in0(N__17762),
            .in1(N__17542),
            .in2(N__17319),
            .in3(N__17590),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_8_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_8_6_6 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_8_6_6  (
            .in0(N__14396),
            .in1(N__16586),
            .in2(N__16634),
            .in3(N__17262),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_6_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_8_6_7  (
            .in0(N__14771),
            .in1(N__16519),
            .in2(N__14755),
            .in3(N__17432),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0  (
            .in0(N__20624),
            .in1(N__21376),
            .in2(N__21277),
            .in3(N__21135),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__18079),
            .in2(_gnd_net_),
            .in3(N__21032),
            .lcout(\Lab_UT.bu_rx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_8_7_2  (
            .in0(N__18119),
            .in1(N__17825),
            .in2(N__18087),
            .in3(N__14713),
            .lcout(\Lab_UT.dictrl.dicLdAMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22305),
            .ce(),
            .sr(N__20943));
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_LC_8_7_3  (
            .in0(N__17826),
            .in1(N__18159),
            .in2(N__14824),
            .in3(N__18083),
            .lcout(\Lab_UT.dictrl.dicRun_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22305),
            .ce(),
            .sr(N__20943));
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6  (
            .in0(N__21255),
            .in1(N__21375),
            .in2(_gnd_net_),
            .in3(N__14712),
            .lcout(\Lab_UT.LdAMones ),
            .ltout(\Lab_UT.LdAMones_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7  (
            .in0(N__14790),
            .in1(N__14808),
            .in2(N__14692),
            .in3(N__18463),
            .lcout(\Lab_UT.loadalarm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_8_8_0 .LUT_INIT=16'b0101010001010111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_LC_8_8_0  (
            .in0(N__19137),
            .in1(N__19267),
            .in2(N__18700),
            .in3(N__15087),
            .lcout(\Lab_UT.dictrl.state_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__18530),
            .sr(N__20937));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_8_8_1 .LUT_INIT=16'b0000000111111101;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_LC_8_8_1  (
            .in0(N__15088),
            .in1(N__18699),
            .in2(N__19275),
            .in3(N__19138),
            .lcout(\Lab_UT.dictrl.state_ret_2_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__18530),
            .sr(N__20937));
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_8_8_3 .LUT_INIT=16'b0000000111111101;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_ess_LC_8_8_3  (
            .in0(N__14872),
            .in1(N__19054),
            .in2(N__19276),
            .in3(N__14848),
            .lcout(\Lab_UT.dictrl.state_i_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__18530),
            .sr(N__20937));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_8_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__18486),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(\Lab_UT.dictrl.m19_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_esr_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_esr_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_esr_LC_8_8_5 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_esr_LC_8_8_5  (
            .in0(N__19266),
            .in1(N__18886),
            .in2(N__18745),
            .in3(N__18158),
            .lcout(\Lab_UT.dictrl.next_state66_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__18530),
            .sr(N__20937));
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_8_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_8_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_RNICG571_LC_8_8_6  (
            .in0(N__14820),
            .in1(N__21226),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\Lab_UT.LdASones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0  (
            .in0(N__15007),
            .in1(N__15046),
            .in2(N__14973),
            .in3(N__18814),
            .lcout(\Lab_UT.next_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1  (
            .in0(N__18817),
            .in1(N__14972),
            .in2(N__15055),
            .in3(N__15010),
            .lcout(\Lab_UT.dictrl.state_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2  (
            .in0(N__15008),
            .in1(N__15047),
            .in2(N__14974),
            .in3(N__18815),
            .lcout(\Lab_UT.dictrl.state_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3  (
            .in0(N__18816),
            .in1(N__14971),
            .in2(N__15054),
            .in3(N__15009),
            .lcout(\Lab_UT.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4  (
            .in0(N__21225),
            .in1(N__20582),
            .in2(N__18559),
            .in3(N__21359),
            .lcout(\Lab_UT.LdAStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5  (
            .in0(N__18879),
            .in1(N__18733),
            .in2(_gnd_net_),
            .in3(N__19227),
            .lcout(\Lab_UT.state_i_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__19226),
            .in2(N__18740),
            .in3(N__18878),
            .lcout(\Lab_UT.dictrl.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7  (
            .in0(N__14867),
            .in1(N__14844),
            .in2(N__19071),
            .in3(N__19228),
            .lcout(Lab_UT_dictrl_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(N__18538),
            .sr(N__20944));
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0  (
            .in0(N__19246),
            .in1(N__14943),
            .in2(N__14932),
            .in3(N__18560),
            .lcout(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_8_10_1  (
            .in0(N__18562),
            .in1(N__19051),
            .in2(N__14871),
            .in3(N__14944),
            .lcout(\Lab_UT.dictrl.next_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22281),
            .ce(N__19331),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2  (
            .in0(N__14904),
            .in1(N__14892),
            .in2(N__15031),
            .in3(N__20613),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_20_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3  (
            .in0(N__18561),
            .in1(N__19049),
            .in2(N__14923),
            .in3(N__14920),
            .lcout(),
            .ltout(\Lab_UT.next_state_1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \Lab_UT.didp.g0_0_LC_8_10_4  (
            .in0(N__18124),
            .in1(N__14914),
            .in2(N__14908),
            .in3(N__17809),
            .lcout(\Lab_UT.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6  (
            .in0(N__14905),
            .in1(N__14893),
            .in2(N__14884),
            .in3(N__20614),
            .lcout(\Lab_UT.dictrl.N_20 ),
            .ltout(\Lab_UT.dictrl.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7  (
            .in0(N__19244),
            .in1(N__14843),
            .in2(N__14827),
            .in3(N__19050),
            .lcout(\Lab_UT.next_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_8_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_8_11_1 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_8_11_1  (
            .in0(N__20310),
            .in1(N__19827),
            .in2(N__20185),
            .in3(N__20030),
            .lcout(N_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_8_11_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_8_11_2  (
            .in0(N__19209),
            .in1(N__18840),
            .in2(N__19294),
            .in3(N__15064),
            .lcout(\Lab_UT.dictrl.G_14_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__18487),
            .in2(_gnd_net_),
            .in3(N__21143),
            .lcout(\Lab_UT.dictrl.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_8_11_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_8_11_4  (
            .in0(N__19828),
            .in1(N__19894),
            .in2(N__15022),
            .in3(N__21425),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_8_11_5 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_8_11_5  (
            .in0(N__18841),
            .in1(N__20621),
            .in2(N__15013),
            .in3(N__14982),
            .lcout(\Lab_UT.dictrl.G_14_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_8_11_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_8_11_6  (
            .in0(N__19208),
            .in1(N__19061),
            .in2(_gnd_net_),
            .in3(N__18936),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_14_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_8_11_7 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_8_11_7  (
            .in0(N__20616),
            .in1(N__14992),
            .in2(N__14986),
            .in3(N__14983),
            .lcout(\Lab_UT.dictrl.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_12_0 .LUT_INIT=16'b1010101011111101;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_12_0  (
            .in0(N__19816),
            .in1(N__19121),
            .in2(N__19730),
            .in3(N__19869),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1  (
            .in0(N__19713),
            .in1(N__15070),
            .in2(N__14947),
            .in3(N__19590),
            .lcout(\Lab_UT.dictrl.N_60_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_2  (
            .in0(N__19062),
            .in1(N__15226),
            .in2(N__15199),
            .in3(N__19631),
            .lcout(\Lab_UT.dictrl.i8_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3  (
            .in0(N__19122),
            .in1(N__20468),
            .in2(_gnd_net_),
            .in3(N__19817),
            .lcout(),
            .ltout(N_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .LUT_INIT=16'b0101000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4  (
            .in0(N__19063),
            .in1(N__18948),
            .in2(N__15133),
            .in3(N__20622),
            .lcout(\Lab_UT.dictrl.G_6_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_8_12_5 .LUT_INIT=16'b0010011110100111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_5_0_LC_8_12_5  (
            .in0(N__21423),
            .in1(N__19818),
            .in2(N__20038),
            .in3(N__19589),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_8_12_6 .LUT_INIT=16'b1111000001111111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_3_0_LC_8_12_6  (
            .in0(N__15130),
            .in1(N__15114),
            .in2(N__15118),
            .in3(N__21424),
            .lcout(\Lab_UT.dictrl.i9_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_8_12_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_8_12_7  (
            .in0(N__20623),
            .in1(N__19064),
            .in2(N__15661),
            .in3(N__15115),
            .lcout(\Lab_UT.dictrl.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_8_13_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_8_13_0  (
            .in0(N__15103),
            .in1(N__15094),
            .in2(_gnd_net_),
            .in3(N__19090),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_13_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_13_1  (
            .in0(N__15711),
            .in1(N__15765),
            .in2(N__19736),
            .in3(N__15405),
            .lcout(\Lab_UT.dictrl.g0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_13_2 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_13_2  (
            .in0(N__19714),
            .in1(N__19112),
            .in2(N__19921),
            .in3(N__19779),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m22_x1_LC_8_13_4  (
            .in0(N__19454),
            .in1(N__20007),
            .in2(N__15784),
            .in3(N__15710),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m22_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.m22_ns_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15415),
            .in3(N__15248),
            .lcout(\Lab_UT.dictrl.N_72_mux ),
            .ltout(\Lab_UT.dictrl.N_72_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__19868),
            .in2(N__15412),
            .in3(N__19778),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_8_14_0 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_8_14_0  (
            .in0(N__15795),
            .in1(N__19464),
            .in2(N__19545),
            .in3(N__15409),
            .lcout(\Lab_UT.dictrl.g0_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_x1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_x1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_x1_LC_8_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_x1_LC_8_14_1  (
            .in0(N__19513),
            .in1(N__15621),
            .in2(N__15331),
            .in3(N__15299),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15280),
            .in3(N__15277),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_3  (
            .in0(N__15232),
            .in1(N__15268),
            .in2(N__15262),
            .in3(N__21426),
            .lcout(\Lab_UT.dictrl.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_4_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_4_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_4_LC_8_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.m22_4_LC_8_14_4  (
            .in0(N__15647),
            .in1(N__19398),
            .in2(N__15625),
            .in3(N__19363),
            .lcout(\Lab_UT.dictrl.m22Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.g0_5_4_LC_8_14_5  (
            .in0(N__19364),
            .in1(N__15623),
            .in2(N__19405),
            .in3(N__19691),
            .lcout(\Lab_UT.dictrl.g0_5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_8_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_8_14_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_8_14_6  (
            .in0(N__20032),
            .in1(N__21431),
            .in2(N__15799),
            .in3(N__15709),
            .lcout(G_6_0_a6_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_7  (
            .in0(N__19399),
            .in1(N__15622),
            .in2(N__19544),
            .in3(N__15648),
            .lcout(\Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15601),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__15474),
            .sr(N__20973));
    defparam \buart.Z_rx.shifter_7_LC_8_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_8_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15600),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__15474),
            .sr(N__20973));
    defparam \buart.Z_rx.shifter_fast_0_LC_8_15_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_8_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20191),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__15474),
            .sr(N__20973));
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15525),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__15474),
            .sr(N__20973));
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0  (
            .in0(N__15988),
            .in1(N__20739),
            .in2(N__15448),
            .in3(N__15967),
            .lcout(\uu2.un3_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_9_1_1  (
            .in0(N__15969),
            .in1(N__15993),
            .in2(N__21952),
            .in3(N__20741),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15853),
            .sr(N__15841));
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2  (
            .in0(N__16012),
            .in1(N__15866),
            .in2(_gnd_net_),
            .in3(N__21946),
            .lcout(),
            .ltout(\uu2.un3_w_addr_user_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.w_addr_user_RNIINVH_4_LC_9_1_3  (
            .in0(N__16048),
            .in1(N__16189),
            .in2(N__16162),
            .in3(N__16159),
            .lcout(\uu2.un3_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_4  (
            .in0(N__15989),
            .in1(N__21903),
            .in2(_gnd_net_),
            .in3(N__16137),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_9_1_5  (
            .in0(N__16049),
            .in1(N__15915),
            .in2(N__16018),
            .in3(N__15903),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15853),
            .sr(N__15841));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_6 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_6  (
            .in0(N__20740),
            .in1(N__21947),
            .in2(N__15994),
            .in3(N__15968),
            .lcout(\uu2.un404_ci ),
            .ltout(\uu2.un404_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_9_1_7  (
            .in0(N__15867),
            .in1(N__15902),
            .in2(N__15880),
            .in3(N__15877),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15853),
            .sr(N__15841));
    defparam \uu2.bitmap_290_LC_9_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_9_2_0 .LUT_INIT=16'b0001001000100111;
    LogicCell40 \uu2.bitmap_290_LC_9_2_0  (
            .in0(N__16557),
            .in1(N__16379),
            .in2(N__17372),
            .in3(N__16416),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_194_LC_9_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_9_2_1 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \uu2.bitmap_194_LC_9_2_1  (
            .in0(N__16415),
            .in1(N__17359),
            .in2(N__16388),
            .in3(N__16556),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_66_LC_9_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_9_2_2 .LUT_INIT=16'b0001010000110101;
    LogicCell40 \uu2.bitmap_66_LC_9_2_2  (
            .in0(N__16559),
            .in1(N__16383),
            .in2(N__17373),
            .in3(N__16418),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_RNIPDM31_66_LC_9_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPDM31_66_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPDM31_66_LC_9_2_3 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \uu2.bitmap_RNIPDM31_66_LC_9_2_3  (
            .in0(N__15811),
            .in1(N__16309),
            .in2(N__16264),
            .in3(N__15805),
            .lcout(\uu2.bitmap_pmux_20_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_9_2_4 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_9_2_4 .LUT_INIT=16'b0001011000110110;
    LogicCell40 \uu2.bitmap_162_LC_9_2_4  (
            .in0(N__16555),
            .in1(N__16375),
            .in2(N__17371),
            .in3(N__16414),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_34_LC_9_2_5 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_9_2_5 .LUT_INIT=16'b1101111101111001;
    LogicCell40 \uu2.bitmap_34_LC_9_2_5  (
            .in0(N__16417),
            .in1(N__17363),
            .in2(N__16389),
            .in3(N__16558),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_RNIP2JO1_34_LC_9_2_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIP2JO1_34_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIP2JO1_34_LC_9_2_6 .LUT_INIT=16'b0000111111001010;
    LogicCell40 \uu2.bitmap_RNIP2JO1_34_LC_9_2_6  (
            .in0(N__16492),
            .in1(N__16486),
            .in2(N__16480),
            .in3(N__16463),
            .lcout(\uu2.bitmap_RNIP2JO1Z0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_69_LC_9_2_7 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_9_2_7 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \uu2.bitmap_69_LC_9_2_7  (
            .in0(N__16419),
            .in1(N__17367),
            .in2(N__16390),
            .in3(N__16560),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20906));
    defparam \uu2.bitmap_314_LC_9_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_9_3_0 .LUT_INIT=16'b0000011000011101;
    LogicCell40 \uu2.bitmap_314_LC_9_3_0  (
            .in0(N__16803),
            .in1(N__16840),
            .in2(N__16883),
            .in3(N__16908),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20904));
    defparam \uu2.bitmap_218_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_9_3_1 .LUT_INIT=16'b0001000000010101;
    LogicCell40 \uu2.bitmap_218_LC_9_3_1  (
            .in0(N__16907),
            .in1(N__16870),
            .in2(N__16845),
            .in3(N__16802),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20904));
    defparam \uu2.bitmap_90_LC_9_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_9_3_2 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \uu2.bitmap_90_LC_9_3_2  (
            .in0(N__16805),
            .in1(N__16844),
            .in2(N__16884),
            .in3(N__16910),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20904));
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \uu2.bitmap_RNIJ4K41_90_LC_9_3_3  (
            .in0(N__16310),
            .in1(N__16270),
            .in2(N__16250),
            .in3(N__16204),
            .lcout(\uu2.bitmap_pmux_19_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_9_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_9_3_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_186_LC_9_3_4  (
            .in0(N__16801),
            .in1(N__16836),
            .in2(N__16882),
            .in3(N__16906),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20904));
    defparam \uu2.bitmap_58_LC_9_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_9_3_5 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_58_LC_9_3_5  (
            .in0(N__16909),
            .in1(N__16874),
            .in2(N__16846),
            .in3(N__16804),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20904));
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNIM5E21_314_LC_9_3_7  (
            .in0(N__16779),
            .in1(N__16765),
            .in2(_gnd_net_),
            .in3(N__16681),
            .lcout(\uu2.bitmap_RNIM5E21Z0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIKGSI_58_LC_9_4_6  (
            .in0(N__16713),
            .in1(N__16693),
            .in2(_gnd_net_),
            .in3(N__16687),
            .lcout(\uu2.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_9_4_7  (
            .in0(N__17968),
            .in1(N__17530),
            .in2(N__18011),
            .in3(N__17176),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22334),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI62AM_1_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__16675),
            .in2(_gnd_net_),
            .in3(N__17869),
            .lcout(\Lab_UT.didp.un1_dicLdStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_9_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_9_5_1  (
            .in0(N__17518),
            .in1(N__16624),
            .in2(_gnd_net_),
            .in3(N__16591),
            .lcout(\Lab_UT.min1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_5_3 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_5_3  (
            .in0(N__17108),
            .in1(N__20341),
            .in2(N__16528),
            .in3(N__17433),
            .lcout(\Lab_UT.didp.countrce4.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4  (
            .in0(N__17002),
            .in1(N__17231),
            .in2(_gnd_net_),
            .in3(N__17933),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5  (
            .in0(N__16941),
            .in1(N__20524),
            .in2(N__17533),
            .in3(N__17175),
            .lcout(\Lab_UT.didp.countrce3.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__17727),
            .in2(_gnd_net_),
            .in3(N__17582),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_5_7 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_5_7  (
            .in0(N__17639),
            .in1(N__20340),
            .in2(N__17524),
            .in3(N__17269),
            .lcout(\Lab_UT.didp.countrce1.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_9_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_9_6_2  (
            .in0(N__17499),
            .in1(N__17430),
            .in2(_gnd_net_),
            .in3(N__17401),
            .lcout(\Lab_UT.min1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_9_6_3  (
            .in0(N__17746),
            .in1(N__17329),
            .in2(N__17323),
            .in3(N__17270),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_6_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_6_4  (
            .in0(N__17000),
            .in1(N__17236),
            .in2(N__17187),
            .in3(N__17930),
            .lcout(\Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_9_6_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_9_6_5  (
            .in0(N__17117),
            .in1(N__20516),
            .in2(N__17059),
            .in3(N__17040),
            .lcout(\Lab_UT.didp.countrce4.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_6 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_6  (
            .in0(N__17001),
            .in1(N__20200),
            .in2(N__16953),
            .in3(N__17931),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_6_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_9_6_7  (
            .in0(N__17932),
            .in1(N__18012),
            .in2(N__17971),
            .in3(N__17964),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_9_7_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_esr_LC_9_7_0  (
            .in0(N__18169),
            .in1(N__17827),
            .in2(N__18861),
            .in3(N__18120),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__18526),
            .sr(N__20946));
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_9_7_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_9_7_1 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_ess_LC_9_7_1  (
            .in0(N__18121),
            .in1(N__18857),
            .in2(N__17835),
            .in3(N__18170),
            .lcout(\Lab_UT.LdSones_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__18526),
            .sr(N__20946));
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_7_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_7_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_LC_9_7_2  (
            .in0(N__18171),
            .in1(N__17831),
            .in2(N__18862),
            .in3(N__18122),
            .lcout(\Lab_UT.state_ret_8_ess ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__18526),
            .sr(N__20946));
    defparam \Lab_UT.didp.state_ret_1_esr_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.state_ret_1_esr_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.state_ret_1_esr_LC_9_7_3 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \Lab_UT.didp.state_ret_1_esr_LC_9_7_3  (
            .in0(N__18123),
            .in1(_gnd_net_),
            .in2(N__17836),
            .in3(N__18172),
            .lcout(\Lab_UT.didp.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__18526),
            .sr(N__20946));
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_9_7_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \Lab_UT.didp.ce_RNIFQ9K_0_LC_9_7_4  (
            .in0(N__17779),
            .in1(N__17770),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.un1_dicLdSones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_7_7 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_7_7  (
            .in0(N__17726),
            .in1(N__20186),
            .in2(N__17638),
            .in3(N__17589),
            .lcout(\Lab_UT.didp.countrce1.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_9_8_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_9_8_0  (
            .in0(N__18495),
            .in1(N__21486),
            .in2(_gnd_net_),
            .in3(N__18670),
            .lcout(\Lab_UT.next_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_9_8_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI81O17_2_LC_9_8_1  (
            .in0(N__19259),
            .in1(N__21307),
            .in2(N__18597),
            .in3(N__21229),
            .lcout(\Lab_UT.dictrl.g0_1_mb_rn_0 ),
            .ltout(\Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_9_8_2 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_2_LC_9_8_2  (
            .in0(N__18496),
            .in1(_gnd_net_),
            .in2(N__18664),
            .in3(N__21487),
            .lcout(\Lab_UT.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22306),
            .ce(N__18537),
            .sr(N__20940));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_9_8_3 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_9_8_3  (
            .in0(N__21108),
            .in1(N__18657),
            .in2(N__18630),
            .in3(N__21230),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_9_8_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_9_8_4 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__18593),
            .in2(N__18565),
            .in3(N__19263),
            .lcout(\Lab_UT.dictrl.state_i_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22306),
            .ce(N__18537),
            .sr(N__20940));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_9_8_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_9_8_5  (
            .in0(N__21107),
            .in1(_gnd_net_),
            .in2(N__19274),
            .in3(N__21228),
            .lcout(\Lab_UT.dictrl.g0_1_mb_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_9_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__18482),
            .in2(_gnd_net_),
            .in3(N__21106),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un15_loadalarm_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_9_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_9_8_7 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_9_8_7  (
            .in0(N__18920),
            .in1(N__21227),
            .in2(N__18466),
            .in3(N__20583),
            .lcout(\Lab_UT.dictrl.loadalarm_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_9_9_2  (
            .in0(N__18457),
            .in1(N__18216),
            .in2(_gnd_net_),
            .in3(N__18370),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22297),
            .ce(),
            .sr(N__20947));
    defparam \Lab_UT.dictrl.state_ret_9_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_LC_9_9_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_9_LC_9_9_4 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_LC_9_9_4  (
            .in0(N__18153),
            .in1(N__18118),
            .in2(N__18088),
            .in3(N__18935),
            .lcout(\Lab_UT.dicLdSones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22297),
            .ce(),
            .sr(N__20947));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__21250),
            .in2(_gnd_net_),
            .in3(N__21373),
            .lcout(\Lab_UT.dictrl.m34_0 ),
            .ltout(\Lab_UT.dictrl.m34_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_9_10_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m35_LC_9_10_2  (
            .in0(N__18801),
            .in1(N__18777),
            .in2(N__18889),
            .in3(N__21141),
            .lcout(\Lab_UT.dictrl.next_state_1_3 ),
            .ltout(\Lab_UT.dictrl.next_state_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_9_10_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__18726),
            .in2(N__18865),
            .in3(N__19231),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_9_10_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_9_10_4  (
            .in0(N__19229),
            .in1(N__19030),
            .in2(_gnd_net_),
            .in3(N__21139),
            .lcout(\Lab_UT.dictrl.N_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_9_10_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_9_10_5  (
            .in0(N__21140),
            .in1(N__19230),
            .in2(_gnd_net_),
            .in3(N__19034),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_9_10_6 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_9_10_6  (
            .in0(N__21374),
            .in1(N__18829),
            .in2(N__18820),
            .in3(N__19555),
            .lcout(\Lab_UT.dictrl.N_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_3_LC_9_10_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_9_10_7  (
            .in0(N__21142),
            .in1(N__18802),
            .in2(N__18787),
            .in3(N__18778),
            .lcout(\Lab_UT.dictrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22289),
            .ce(N__19327),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_2  (
            .in0(N__20532),
            .in1(_gnd_net_),
            .in2(N__18970),
            .in3(N__21418),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__18695),
            .in2(N__19345),
            .in3(N__18895),
            .lcout(\Lab_UT.dictrl.next_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(N__19341),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6  (
            .in0(N__19290),
            .in1(N__19264),
            .in2(_gnd_net_),
            .in3(N__21417),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7  (
            .in0(N__19265),
            .in1(N__18965),
            .in2(N__19141),
            .in3(N__20533),
            .lcout(\Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m7_0_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m7_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m7_0_LC_9_12_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.m7_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__19123),
            .in2(_gnd_net_),
            .in3(N__19826),
            .lcout(\Lab_UT.dictrl.N_8_0 ),
            .ltout(\Lab_UT.dictrl.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_12_1 .LUT_INIT=16'b1100110010101111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_12_1  (
            .in0(N__20498),
            .in1(N__20352),
            .in2(N__19096),
            .in3(N__20618),
            .lcout(\Lab_UT.dictrl.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_2 .LUT_INIT=16'b0111010101110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_2  (
            .in0(N__20617),
            .in1(N__18937),
            .in2(N__19072),
            .in3(N__21416),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_6_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .LUT_INIT=16'b0011010000000100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3  (
            .in0(N__20359),
            .in1(N__19068),
            .in2(N__19093),
            .in3(N__19930),
            .lcout(\Lab_UT.dictrl.G_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_5 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_5  (
            .in0(N__19084),
            .in1(N__19078),
            .in2(N__20517),
            .in3(N__20620),
            .lcout(),
            .ltout(\Lab_UT.dictrl.i8_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_12_6 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_12_6  (
            .in0(N__19069),
            .in1(N__18969),
            .in2(N__18952),
            .in3(N__18938),
            .lcout(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_7  (
            .in0(N__20358),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__20619),
            .lcout(\Lab_UT.dictrl.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m14_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m14_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m14_LC_9_13_1 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \Lab_UT.dictrl.m14_LC_9_13_1  (
            .in0(N__19824),
            .in1(N__20494),
            .in2(_gnd_net_),
            .in3(N__19597),
            .lcout(\Lab_UT.dictrl.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_13_2 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_13_2  (
            .in0(N__20302),
            .in1(N__19825),
            .in2(N__20198),
            .in3(N__20031),
            .lcout(G_6_0_a6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_9_13_6 .LUT_INIT=16'b1111101101010001;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_9_13_6  (
            .in0(N__19918),
            .in1(N__19823),
            .in2(N__19737),
            .in3(N__19627),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_9_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_9_13_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__19606),
            .in2(N__19600),
            .in3(N__19596),
            .lcout(\Lab_UT.dictrl.N_59_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_9_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_9_14_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_9_14_0  (
            .in0(N__19546),
            .in1(N__19512),
            .in2(_gnd_net_),
            .in3(N__19498),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_9_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_9_14_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_9_14_1  (
            .in0(N__19477),
            .in1(N__19465),
            .in2(N__19408),
            .in3(N__19404),
            .lcout(\Lab_UT.dictrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_9_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_9_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_9_14_3  (
            .in0(N__19378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19372),
            .lcout(\Lab_UT.dictrl.g0_6_3 ),
            .ltout(\Lab_UT.dictrl.g0_6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_9_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_9_14_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_9_14_4  (
            .in0(N__21456),
            .in1(N__21466),
            .in2(N__21490),
            .in3(N__21442),
            .lcout(\Lab_UT.dictrl.N_57_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_9_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_9_14_6 .LUT_INIT=16'b0101111100110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_8_LC_9_14_6  (
            .in0(N__21472),
            .in1(N__21465),
            .in2(N__21457),
            .in3(N__21441),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_9_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_9_14_7 .LUT_INIT=16'b0011111101110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_4_LC_9_14_7  (
            .in0(N__21303),
            .in1(N__21283),
            .in2(N__21172),
            .in3(N__21153),
            .lcout(\Lab_UT.dictrl.G_25_i_a5_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .LUT_INIT=16'b1111100111111100;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_11_1_0  (
            .in0(N__21517),
            .in1(N__21556),
            .in2(N__21714),
            .in3(N__21578),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(N__20974));
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_11_1_1  (
            .in0(N__21577),
            .in1(N__21698),
            .in2(_gnd_net_),
            .in3(N__21516),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(N__20974));
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_11_1_2  (
            .in0(N__21595),
            .in1(N__21496),
            .in2(N__21715),
            .in3(N__21580),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(N__20974));
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .LUT_INIT=16'b0000000010010110;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_11_1_3  (
            .in0(N__21579),
            .in1(N__21721),
            .in2(N__21538),
            .in3(N__21702),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(N__20974));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5  (
            .in0(N__20742),
            .in1(N__21917),
            .in2(_gnd_net_),
            .in3(N__20704),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7  (
            .in0(N__21951),
            .in1(N__21918),
            .in2(_gnd_net_),
            .in3(N__21799),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0  (
            .in0(N__21514),
            .in1(N__21554),
            .in2(_gnd_net_),
            .in3(N__21575),
            .lcout(\buart.Z_tx.un1_bitcount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__22027),
            .in2(_gnd_net_),
            .in3(N__22011),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22347),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_2_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__21678),
            .in2(_gnd_net_),
            .in3(N__21576),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22010),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22347),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__21594),
            .in2(_gnd_net_),
            .in3(N__21513),
            .lcout(),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6  (
            .in0(N__21533),
            .in1(N__21553),
            .in2(N__21583),
            .in3(N__21967),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7  (
            .in0(N__21555),
            .in1(N__21534),
            .in2(N__21520),
            .in3(N__21515),
            .lcout(\buart.Z_tx.un1_bitcount_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__22026),
            .in2(N__22012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21991),
            .in3(N__22372),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__22350),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2  (
            .in0(N__21969),
            .in1(N__22036),
            .in2(_gnd_net_),
            .in3(N__22369),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__22350),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22063),
            .in3(N__22366),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__22350),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4  (
            .in0(N__21970),
            .in1(_gnd_net_),
            .in2(N__22075),
            .in3(N__22363),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__22350),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5  (
            .in0(N__22050),
            .in1(N__21968),
            .in2(_gnd_net_),
            .in3(N__22360),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22350),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6  (
            .in0(N__22071),
            .in1(N__22059),
            .in2(N__22051),
            .in3(N__22035),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7  (
            .in0(N__22025),
            .in1(N__22006),
            .in2(N__21990),
            .in3(N__21976),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
