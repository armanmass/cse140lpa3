// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 19 2019 22:38:34

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__23331;
    wire N__23330;
    wire N__23329;
    wire N__23322;
    wire N__23321;
    wire N__23320;
    wire N__23313;
    wire N__23312;
    wire N__23311;
    wire N__23304;
    wire N__23303;
    wire N__23302;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23277;
    wire N__23276;
    wire N__23275;
    wire N__23268;
    wire N__23267;
    wire N__23266;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23209;
    wire N__23206;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23199;
    wire N__23198;
    wire N__23197;
    wire N__23196;
    wire N__23195;
    wire N__23194;
    wire N__23193;
    wire N__23192;
    wire N__23189;
    wire N__23182;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23170;
    wire N__23167;
    wire N__23160;
    wire N__23155;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23130;
    wire N__23125;
    wire N__23122;
    wire N__23117;
    wire N__23108;
    wire N__23105;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23086;
    wire N__23085;
    wire N__23084;
    wire N__23083;
    wire N__23080;
    wire N__23079;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23042;
    wire N__23035;
    wire N__23034;
    wire N__23033;
    wire N__23030;
    wire N__23025;
    wire N__23022;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22994;
    wire N__22989;
    wire N__22976;
    wire N__22975;
    wire N__22974;
    wire N__22973;
    wire N__22972;
    wire N__22971;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22965;
    wire N__22962;
    wire N__22961;
    wire N__22960;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22941;
    wire N__22938;
    wire N__22933;
    wire N__22930;
    wire N__22925;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22886;
    wire N__22877;
    wire N__22876;
    wire N__22875;
    wire N__22872;
    wire N__22871;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22863;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22824;
    wire N__22821;
    wire N__22814;
    wire N__22809;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22793;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22769;
    wire N__22768;
    wire N__22767;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22760;
    wire N__22759;
    wire N__22756;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22748;
    wire N__22747;
    wire N__22744;
    wire N__22743;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22736;
    wire N__22733;
    wire N__22728;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22702;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22672;
    wire N__22665;
    wire N__22660;
    wire N__22655;
    wire N__22652;
    wire N__22647;
    wire N__22642;
    wire N__22635;
    wire N__22630;
    wire N__22627;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22599;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22559;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22546;
    wire N__22545;
    wire N__22544;
    wire N__22541;
    wire N__22536;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22528;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22520;
    wire N__22513;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22499;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22483;
    wire N__22476;
    wire N__22471;
    wire N__22460;
    wire N__22459;
    wire N__22458;
    wire N__22457;
    wire N__22456;
    wire N__22455;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22436;
    wire N__22435;
    wire N__22434;
    wire N__22431;
    wire N__22430;
    wire N__22427;
    wire N__22420;
    wire N__22419;
    wire N__22416;
    wire N__22409;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22380;
    wire N__22375;
    wire N__22372;
    wire N__22361;
    wire N__22360;
    wire N__22359;
    wire N__22358;
    wire N__22357;
    wire N__22356;
    wire N__22355;
    wire N__22354;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22350;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22346;
    wire N__22345;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22337;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22330;
    wire N__22329;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22317;
    wire N__22316;
    wire N__22315;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22311;
    wire N__22310;
    wire N__22309;
    wire N__22308;
    wire N__22307;
    wire N__22306;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22301;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22275;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22075;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22070;
    wire N__22069;
    wire N__22068;
    wire N__22067;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22039;
    wire N__22038;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22014;
    wire N__22013;
    wire N__22012;
    wire N__22011;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22007;
    wire N__22006;
    wire N__22005;
    wire N__22004;
    wire N__22003;
    wire N__22002;
    wire N__22001;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21973;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21940;
    wire N__21939;
    wire N__21938;
    wire N__21935;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21785;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21754;
    wire N__21753;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21741;
    wire N__21740;
    wire N__21739;
    wire N__21738;
    wire N__21729;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21694;
    wire N__21693;
    wire N__21686;
    wire N__21679;
    wire N__21674;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21623;
    wire N__21620;
    wire N__21619;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21598;
    wire N__21591;
    wire N__21588;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21564;
    wire N__21561;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21535;
    wire N__21534;
    wire N__21531;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21508;
    wire N__21503;
    wire N__21500;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21456;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21435;
    wire N__21434;
    wire N__21433;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21411;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21392;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21377;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21373;
    wire N__21370;
    wire N__21369;
    wire N__21366;
    wire N__21365;
    wire N__21364;
    wire N__21363;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21310;
    wire N__21307;
    wire N__21296;
    wire N__21281;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21203;
    wire N__21202;
    wire N__21199;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21182;
    wire N__21179;
    wire N__21174;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21147;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21125;
    wire N__21124;
    wire N__21123;
    wire N__21118;
    wire N__21115;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21105;
    wire N__21100;
    wire N__21095;
    wire N__21092;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21068;
    wire N__21067;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21051;
    wire N__21048;
    wire N__21043;
    wire N__21036;
    wire N__21033;
    wire N__21028;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21010;
    wire N__21007;
    wire N__21002;
    wire N__20995;
    wire N__20988;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20954;
    wire N__20953;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20949;
    wire N__20944;
    wire N__20943;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20853;
    wire N__20852;
    wire N__20851;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20833;
    wire N__20830;
    wire N__20829;
    wire N__20828;
    wire N__20825;
    wire N__20818;
    wire N__20817;
    wire N__20812;
    wire N__20811;
    wire N__20808;
    wire N__20801;
    wire N__20800;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20795;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20764;
    wire N__20761;
    wire N__20756;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20728;
    wire N__20727;
    wire N__20726;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20698;
    wire N__20695;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20659;
    wire N__20658;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20654;
    wire N__20651;
    wire N__20650;
    wire N__20649;
    wire N__20646;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20628;
    wire N__20623;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20606;
    wire N__20605;
    wire N__20604;
    wire N__20603;
    wire N__20602;
    wire N__20601;
    wire N__20598;
    wire N__20591;
    wire N__20586;
    wire N__20583;
    wire N__20578;
    wire N__20573;
    wire N__20570;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20548;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20492;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20482;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20464;
    wire N__20463;
    wire N__20462;
    wire N__20461;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20446;
    wire N__20441;
    wire N__20436;
    wire N__20433;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20391;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20373;
    wire N__20368;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20335;
    wire N__20320;
    wire N__20317;
    wire N__20316;
    wire N__20313;
    wire N__20312;
    wire N__20311;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20293;
    wire N__20290;
    wire N__20285;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20273;
    wire N__20272;
    wire N__20269;
    wire N__20268;
    wire N__20265;
    wire N__20264;
    wire N__20261;
    wire N__20246;
    wire N__20243;
    wire N__20242;
    wire N__20241;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20229;
    wire N__20226;
    wire N__20219;
    wire N__20218;
    wire N__20217;
    wire N__20216;
    wire N__20215;
    wire N__20214;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20194;
    wire N__20185;
    wire N__20184;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20174;
    wire N__20173;
    wire N__20172;
    wire N__20169;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20147;
    wire N__20146;
    wire N__20145;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20131;
    wire N__20124;
    wire N__20123;
    wire N__20120;
    wire N__20115;
    wire N__20112;
    wire N__20111;
    wire N__20110;
    wire N__20109;
    wire N__20108;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20093;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20069;
    wire N__20066;
    wire N__20065;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20054;
    wire N__20053;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20030;
    wire N__20025;
    wire N__20024;
    wire N__20023;
    wire N__20022;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__19999;
    wire N__19996;
    wire N__19989;
    wire N__19982;
    wire N__19981;
    wire N__19980;
    wire N__19979;
    wire N__19978;
    wire N__19977;
    wire N__19976;
    wire N__19975;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19963;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19937;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19909;
    wire N__19908;
    wire N__19907;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19873;
    wire N__19872;
    wire N__19871;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19856;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19833;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19805;
    wire N__19800;
    wire N__19797;
    wire N__19792;
    wire N__19789;
    wire N__19784;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19742;
    wire N__19735;
    wire N__19730;
    wire N__19723;
    wire N__19712;
    wire N__19709;
    wire N__19708;
    wire N__19707;
    wire N__19700;
    wire N__19699;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19678;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19600;
    wire N__19599;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19577;
    wire N__19572;
    wire N__19565;
    wire N__19556;
    wire N__19553;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19543;
    wire N__19542;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19527;
    wire N__19520;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19504;
    wire N__19503;
    wire N__19500;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19450;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19438;
    wire N__19433;
    wire N__19424;
    wire N__19423;
    wire N__19420;
    wire N__19419;
    wire N__19418;
    wire N__19415;
    wire N__19414;
    wire N__19413;
    wire N__19412;
    wire N__19411;
    wire N__19408;
    wire N__19407;
    wire N__19406;
    wire N__19403;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19352;
    wire N__19347;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19326;
    wire N__19325;
    wire N__19324;
    wire N__19323;
    wire N__19322;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19306;
    wire N__19301;
    wire N__19294;
    wire N__19291;
    wire N__19282;
    wire N__19279;
    wire N__19270;
    wire N__19265;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19234;
    wire N__19229;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19207;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19175;
    wire N__19172;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19160;
    wire N__19157;
    wire N__19152;
    wire N__19149;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19120;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19094;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19018;
    wire N__19017;
    wire N__19014;
    wire N__19013;
    wire N__19012;
    wire N__19011;
    wire N__19006;
    wire N__19005;
    wire N__19002;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18967;
    wire N__18962;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18941;
    wire N__18940;
    wire N__18939;
    wire N__18938;
    wire N__18935;
    wire N__18934;
    wire N__18931;
    wire N__18926;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18876;
    wire N__18875;
    wire N__18872;
    wire N__18867;
    wire N__18864;
    wire N__18859;
    wire N__18856;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18831;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18799;
    wire N__18796;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18770;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18705;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18676;
    wire N__18671;
    wire N__18670;
    wire N__18669;
    wire N__18666;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18547;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18542;
    wire N__18527;
    wire N__18526;
    wire N__18525;
    wire N__18524;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18497;
    wire N__18496;
    wire N__18495;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18481;
    wire N__18466;
    wire N__18465;
    wire N__18464;
    wire N__18463;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18448;
    wire N__18445;
    wire N__18440;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18415;
    wire N__18414;
    wire N__18413;
    wire N__18398;
    wire N__18397;
    wire N__18396;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18371;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18367;
    wire N__18366;
    wire N__18365;
    wire N__18364;
    wire N__18349;
    wire N__18348;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18331;
    wire N__18328;
    wire N__18323;
    wire N__18320;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18292;
    wire N__18289;
    wire N__18288;
    wire N__18285;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18250;
    wire N__18245;
    wire N__18242;
    wire N__18241;
    wire N__18238;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18232;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18200;
    wire N__18197;
    wire N__18196;
    wire N__18191;
    wire N__18188;
    wire N__18187;
    wire N__18184;
    wire N__18183;
    wire N__18182;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18165;
    wire N__18160;
    wire N__18157;
    wire N__18146;
    wire N__18145;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18119;
    wire N__18118;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18104;
    wire N__18103;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18091;
    wire N__18088;
    wire N__18081;
    wire N__18076;
    wire N__18073;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18042;
    wire N__18033;
    wire N__18026;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17991;
    wire N__17990;
    wire N__17989;
    wire N__17988;
    wire N__17987;
    wire N__17986;
    wire N__17985;
    wire N__17978;
    wire N__17977;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17952;
    wire N__17947;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17919;
    wire N__17918;
    wire N__17917;
    wire N__17914;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17910;
    wire N__17905;
    wire N__17904;
    wire N__17903;
    wire N__17900;
    wire N__17891;
    wire N__17890;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17866;
    wire N__17865;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17839;
    wire N__17836;
    wire N__17833;
    wire N__17824;
    wire N__17821;
    wire N__17804;
    wire N__17801;
    wire N__17800;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17785;
    wire N__17782;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17764;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17758;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17750;
    wire N__17749;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17728;
    wire N__17723;
    wire N__17718;
    wire N__17715;
    wire N__17710;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17671;
    wire N__17666;
    wire N__17663;
    wire N__17662;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17632;
    wire N__17631;
    wire N__17630;
    wire N__17629;
    wire N__17628;
    wire N__17627;
    wire N__17624;
    wire N__17619;
    wire N__17616;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17557;
    wire N__17552;
    wire N__17551;
    wire N__17548;
    wire N__17547;
    wire N__17546;
    wire N__17545;
    wire N__17542;
    wire N__17541;
    wire N__17538;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17516;
    wire N__17515;
    wire N__17514;
    wire N__17513;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17501;
    wire N__17498;
    wire N__17493;
    wire N__17492;
    wire N__17491;
    wire N__17490;
    wire N__17489;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17485;
    wire N__17484;
    wire N__17477;
    wire N__17476;
    wire N__17473;
    wire N__17468;
    wire N__17459;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17425;
    wire N__17424;
    wire N__17423;
    wire N__17422;
    wire N__17421;
    wire N__17420;
    wire N__17419;
    wire N__17418;
    wire N__17411;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17396;
    wire N__17395;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17389;
    wire N__17388;
    wire N__17387;
    wire N__17382;
    wire N__17379;
    wire N__17374;
    wire N__17369;
    wire N__17366;
    wire N__17359;
    wire N__17354;
    wire N__17351;
    wire N__17344;
    wire N__17333;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17321;
    wire N__17320;
    wire N__17317;
    wire N__17316;
    wire N__17315;
    wire N__17314;
    wire N__17307;
    wire N__17304;
    wire N__17303;
    wire N__17302;
    wire N__17299;
    wire N__17298;
    wire N__17297;
    wire N__17296;
    wire N__17293;
    wire N__17282;
    wire N__17281;
    wire N__17276;
    wire N__17271;
    wire N__17268;
    wire N__17261;
    wire N__17258;
    wire N__17257;
    wire N__17256;
    wire N__17255;
    wire N__17254;
    wire N__17253;
    wire N__17250;
    wire N__17249;
    wire N__17248;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17207;
    wire N__17206;
    wire N__17205;
    wire N__17204;
    wire N__17203;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17189;
    wire N__17186;
    wire N__17181;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17175;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17166;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17147;
    wire N__17144;
    wire N__17139;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17104;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16969;
    wire N__16968;
    wire N__16967;
    wire N__16966;
    wire N__16963;
    wire N__16962;
    wire N__16961;
    wire N__16958;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16950;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16932;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16891;
    wire N__16886;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16861;
    wire N__16860;
    wire N__16859;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16843;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16810;
    wire N__16805;
    wire N__16802;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16790;
    wire N__16787;
    wire N__16786;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16714;
    wire N__16713;
    wire N__16712;
    wire N__16711;
    wire N__16708;
    wire N__16703;
    wire N__16696;
    wire N__16691;
    wire N__16682;
    wire N__16681;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16665;
    wire N__16664;
    wire N__16663;
    wire N__16660;
    wire N__16659;
    wire N__16656;
    wire N__16655;
    wire N__16654;
    wire N__16647;
    wire N__16644;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16594;
    wire N__16593;
    wire N__16592;
    wire N__16591;
    wire N__16584;
    wire N__16579;
    wire N__16578;
    wire N__16577;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16563;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16492;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16483;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16475;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16451;
    wire N__16450;
    wire N__16447;
    wire N__16440;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16424;
    wire N__16415;
    wire N__16414;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16390;
    wire N__16389;
    wire N__16386;
    wire N__16385;
    wire N__16382;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16335;
    wire N__16334;
    wire N__16331;
    wire N__16326;
    wire N__16323;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16305;
    wire N__16302;
    wire N__16301;
    wire N__16300;
    wire N__16299;
    wire N__16294;
    wire N__16293;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16281;
    wire N__16274;
    wire N__16271;
    wire N__16266;
    wire N__16259;
    wire N__16250;
    wire N__16249;
    wire N__16248;
    wire N__16247;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16126;
    wire N__16125;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16110;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16095;
    wire N__16090;
    wire N__16083;
    wire N__16076;
    wire N__16073;
    wire N__16058;
    wire N__16055;
    wire N__16054;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16042;
    wire N__16041;
    wire N__16040;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16028;
    wire N__16025;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16009;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15989;
    wire N__15988;
    wire N__15987;
    wire N__15986;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15974;
    wire N__15969;
    wire N__15962;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15948;
    wire N__15947;
    wire N__15944;
    wire N__15933;
    wire N__15930;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15912;
    wire N__15903;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15881;
    wire N__15876;
    wire N__15873;
    wire N__15860;
    wire N__15859;
    wire N__15858;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15838;
    wire N__15837;
    wire N__15836;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15825;
    wire N__15822;
    wire N__15815;
    wire N__15804;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15778;
    wire N__15775;
    wire N__15770;
    wire N__15755;
    wire N__15754;
    wire N__15749;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15725;
    wire N__15724;
    wire N__15723;
    wire N__15722;
    wire N__15719;
    wire N__15718;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15685;
    wire N__15682;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15671;
    wire N__15668;
    wire N__15659;
    wire N__15658;
    wire N__15657;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15645;
    wire N__15638;
    wire N__15633;
    wire N__15630;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15454;
    wire N__15453;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15441;
    wire N__15440;
    wire N__15437;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15421;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15400;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15376;
    wire N__15373;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15349;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15268;
    wire N__15267;
    wire N__15264;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15252;
    wire N__15249;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15229;
    wire N__15224;
    wire N__15223;
    wire N__15222;
    wire N__15221;
    wire N__15220;
    wire N__15219;
    wire N__15218;
    wire N__15217;
    wire N__15216;
    wire N__15215;
    wire N__15214;
    wire N__15213;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15195;
    wire N__15180;
    wire N__15175;
    wire N__15164;
    wire N__15163;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15159;
    wire N__15158;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15140;
    wire N__15139;
    wire N__15136;
    wire N__15131;
    wire N__15126;
    wire N__15123;
    wire N__15116;
    wire N__15115;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15110;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15086;
    wire N__15083;
    wire N__15076;
    wire N__15067;
    wire N__15064;
    wire N__15059;
    wire N__15054;
    wire N__15047;
    wire N__15046;
    wire N__15043;
    wire N__15042;
    wire N__15037;
    wire N__15034;
    wire N__15033;
    wire N__15032;
    wire N__15029;
    wire N__15028;
    wire N__15027;
    wire N__15026;
    wire N__15025;
    wire N__15024;
    wire N__15023;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15003;
    wire N__14994;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14942;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14908;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14882;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14871;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14859;
    wire N__14856;
    wire N__14849;
    wire N__14846;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14815;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14794;
    wire N__14793;
    wire N__14792;
    wire N__14791;
    wire N__14790;
    wire N__14779;
    wire N__14776;
    wire N__14775;
    wire N__14774;
    wire N__14771;
    wire N__14764;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14718;
    wire N__14715;
    wire N__14714;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14682;
    wire N__14675;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14657;
    wire N__14654;
    wire N__14653;
    wire N__14652;
    wire N__14651;
    wire N__14642;
    wire N__14639;
    wire N__14638;
    wire N__14635;
    wire N__14634;
    wire N__14631;
    wire N__14626;
    wire N__14621;
    wire N__14620;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14594;
    wire N__14591;
    wire N__14590;
    wire N__14589;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14568;
    wire N__14561;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14549;
    wire N__14548;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14498;
    wire N__14497;
    wire N__14496;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14484;
    wire N__14483;
    wire N__14480;
    wire N__14475;
    wire N__14472;
    wire N__14465;
    wire N__14464;
    wire N__14461;
    wire N__14460;
    wire N__14459;
    wire N__14456;
    wire N__14451;
    wire N__14446;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14410;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14384;
    wire N__14381;
    wire N__14374;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14363;
    wire N__14360;
    wire N__14355;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14341;
    wire N__14340;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14306;
    wire N__14305;
    wire N__14302;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14294;
    wire N__14291;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14248;
    wire N__14245;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14223;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14209;
    wire N__14208;
    wire N__14207;
    wire N__14204;
    wire N__14199;
    wire N__14196;
    wire N__14191;
    wire N__14186;
    wire N__14183;
    wire N__14182;
    wire N__14181;
    wire N__14178;
    wire N__14177;
    wire N__14174;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14159;
    wire N__14154;
    wire N__14151;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14123;
    wire N__14122;
    wire N__14121;
    wire N__14120;
    wire N__14119;
    wire N__14112;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14090;
    wire N__14087;
    wire N__14086;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14047;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13948;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13933;
    wire N__13932;
    wire N__13931;
    wire N__13930;
    wire N__13929;
    wire N__13928;
    wire N__13921;
    wire N__13912;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13876;
    wire N__13875;
    wire N__13868;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13846;
    wire N__13845;
    wire N__13844;
    wire N__13843;
    wire N__13842;
    wire N__13837;
    wire N__13828;
    wire N__13823;
    wire N__13820;
    wire N__13819;
    wire N__13818;
    wire N__13817;
    wire N__13814;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13790;
    wire N__13787;
    wire N__13786;
    wire N__13777;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13765;
    wire N__13764;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13739;
    wire N__13738;
    wire N__13737;
    wire N__13734;
    wire N__13729;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13719;
    wire N__13714;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13691;
    wire N__13690;
    wire N__13689;
    wire N__13686;
    wire N__13681;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13655;
    wire N__13652;
    wire N__13651;
    wire N__13650;
    wire N__13647;
    wire N__13642;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13627;
    wire N__13624;
    wire N__13623;
    wire N__13620;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13608;
    wire N__13601;
    wire N__13600;
    wire N__13599;
    wire N__13598;
    wire N__13595;
    wire N__13590;
    wire N__13589;
    wire N__13588;
    wire N__13587;
    wire N__13586;
    wire N__13585;
    wire N__13582;
    wire N__13581;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13560;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13532;
    wire N__13529;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13465;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13448;
    wire N__13443;
    wire N__13438;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13396;
    wire N__13391;
    wire N__13390;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13384;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13364;
    wire N__13361;
    wire N__13360;
    wire N__13359;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13343;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13335;
    wire N__13334;
    wire N__13329;
    wire N__13328;
    wire N__13327;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13290;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13277;
    wire N__13276;
    wire N__13275;
    wire N__13274;
    wire N__13265;
    wire N__13262;
    wire N__13257;
    wire N__13254;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13225;
    wire N__13222;
    wire N__13221;
    wire N__13220;
    wire N__13217;
    wire N__13216;
    wire N__13215;
    wire N__13210;
    wire N__13201;
    wire N__13196;
    wire N__13193;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13181;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13153;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13135;
    wire N__13134;
    wire N__13133;
    wire N__13132;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13120;
    wire N__13115;
    wire N__13110;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13093;
    wire N__13090;
    wire N__13089;
    wire N__13086;
    wire N__13085;
    wire N__13084;
    wire N__13069;
    wire N__13068;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13041;
    wire N__13038;
    wire N__13025;
    wire N__13024;
    wire N__13023;
    wire N__13022;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13014;
    wire N__13013;
    wire N__13010;
    wire N__13009;
    wire N__13006;
    wire N__13005;
    wire N__13004;
    wire N__13001;
    wire N__12986;
    wire N__12981;
    wire N__12976;
    wire N__12971;
    wire N__12970;
    wire N__12969;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12928;
    wire N__12923;
    wire N__12920;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12895;
    wire N__12892;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12867;
    wire N__12864;
    wire N__12859;
    wire N__12854;
    wire N__12853;
    wire N__12852;
    wire N__12851;
    wire N__12850;
    wire N__12845;
    wire N__12840;
    wire N__12837;
    wire N__12830;
    wire N__12829;
    wire N__12828;
    wire N__12827;
    wire N__12824;
    wire N__12823;
    wire N__12816;
    wire N__12811;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12795;
    wire N__12790;
    wire N__12785;
    wire N__12782;
    wire N__12781;
    wire N__12778;
    wire N__12777;
    wire N__12774;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12762;
    wire N__12755;
    wire N__12754;
    wire N__12749;
    wire N__12746;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12729;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12695;
    wire N__12694;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12657;
    wire N__12652;
    wire N__12649;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12613;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12562;
    wire N__12557;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12526;
    wire N__12525;
    wire N__12522;
    wire N__12517;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12482;
    wire N__12481;
    wire N__12480;
    wire N__12477;
    wire N__12472;
    wire N__12467;
    wire N__12464;
    wire N__12463;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12436;
    wire N__12433;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12421;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12295;
    wire N__12290;
    wire N__12287;
    wire N__12286;
    wire N__12281;
    wire N__12278;
    wire N__12277;
    wire N__12274;
    wire N__12269;
    wire N__12266;
    wire N__12265;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12208;
    wire N__12207;
    wire N__12206;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12183;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12149;
    wire N__12148;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12136;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12119;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12100;
    wire N__12097;
    wire N__12092;
    wire N__12091;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__12074;
    wire N__12071;
    wire N__12064;
    wire N__12059;
    wire N__12056;
    wire N__12055;
    wire N__12054;
    wire N__12051;
    wire N__12046;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12031;
    wire N__12028;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12008;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11989;
    wire N__11984;
    wire N__11981;
    wire N__11980;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11965;
    wire N__11960;
    wire N__11959;
    wire N__11956;
    wire N__11955;
    wire N__11948;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11926;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11902;
    wire N__11897;
    wire N__11894;
    wire N__11893;
    wire N__11890;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11858;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11843;
    wire N__11842;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11816;
    wire N__11813;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11774;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11699;
    wire N__11696;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11684;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11579;
    wire N__11574;
    wire N__11571;
    wire N__11564;
    wire N__11555;
    wire N__11548;
    wire N__11547;
    wire N__11544;
    wire N__11541;
    wire N__11536;
    wire N__11527;
    wire N__11524;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11476;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11465;
    wire N__11460;
    wire N__11457;
    wire N__11450;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11438;
    wire N__11431;
    wire N__11426;
    wire N__11423;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11407;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11330;
    wire N__11329;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11308;
    wire N__11305;
    wire N__11300;
    wire N__11297;
    wire N__11292;
    wire N__11287;
    wire N__11282;
    wire N__11273;
    wire N__11270;
    wire N__11269;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11228;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11083;
    wire N__11078;
    wire N__11073;
    wire N__11070;
    wire N__11063;
    wire N__11062;
    wire N__11059;
    wire N__11058;
    wire N__11051;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11036;
    wire N__11035;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11015;
    wire N__11006;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10952;
    wire N__10949;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10917;
    wire N__10916;
    wire N__10915;
    wire N__10912;
    wire N__10903;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10874;
    wire N__10871;
    wire N__10864;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10825;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10807;
    wire N__10802;
    wire N__10799;
    wire N__10798;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10769;
    wire N__10762;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10589;
    wire N__10586;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10548;
    wire N__10545;
    wire N__10544;
    wire N__10539;
    wire N__10534;
    wire N__10531;
    wire N__10526;
    wire N__10517;
    wire N__10514;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10502;
    wire N__10495;
    wire N__10490;
    wire N__10489;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10481;
    wire N__10480;
    wire N__10479;
    wire N__10476;
    wire N__10471;
    wire N__10468;
    wire N__10463;
    wire N__10460;
    wire N__10451;
    wire N__10450;
    wire N__10449;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10430;
    wire N__10427;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10285;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10203;
    wire N__10198;
    wire N__10197;
    wire N__10194;
    wire N__10193;
    wire N__10190;
    wire N__10183;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10143;
    wire N__10138;
    wire N__10133;
    wire N__10132;
    wire N__10127;
    wire N__10126;
    wire N__10125;
    wire N__10122;
    wire N__10117;
    wire N__10112;
    wire N__10111;
    wire N__10110;
    wire N__10109;
    wire N__10108;
    wire N__10105;
    wire N__10100;
    wire N__10095;
    wire N__10092;
    wire N__10087;
    wire N__10082;
    wire N__10079;
    wire N__10078;
    wire N__10077;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10053;
    wire N__10046;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10040;
    wire N__10037;
    wire N__10032;
    wire N__10029;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9996;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9976;
    wire N__9971;
    wire N__9966;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9942;
    wire N__9935;
    wire N__9930;
    wire N__9923;
    wire N__9922;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9904;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9886;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9878;
    wire N__9875;
    wire N__9870;
    wire N__9865;
    wire N__9860;
    wire N__9859;
    wire N__9858;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9812;
    wire N__9809;
    wire N__9808;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9765;
    wire N__9762;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9730;
    wire N__9727;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9696;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9680;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9641;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9616;
    wire N__9607;
    wire N__9602;
    wire N__9599;
    wire N__9590;
    wire N__9587;
    wire N__9578;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9569;
    wire N__9562;
    wire N__9561;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9553;
    wire N__9546;
    wire N__9543;
    wire N__9538;
    wire N__9531;
    wire N__9528;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9473;
    wire N__9472;
    wire N__9471;
    wire N__9470;
    wire N__9461;
    wire N__9458;
    wire N__9457;
    wire N__9456;
    wire N__9453;
    wire N__9448;
    wire N__9445;
    wire N__9440;
    wire N__9439;
    wire N__9438;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9426;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9394;
    wire N__9391;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9373;
    wire N__9364;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9141;
    wire N__9134;
    wire N__9133;
    wire N__9132;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9109;
    wire N__9098;
    wire N__9097;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9000;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8972;
    wire N__8969;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8942;
    wire N__8941;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8924;
    wire N__8923;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8909;
    wire N__8906;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8890;
    wire N__8887;
    wire N__8882;
    wire N__8881;
    wire N__8880;
    wire N__8879;
    wire N__8878;
    wire N__8867;
    wire N__8864;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8854;
    wire N__8851;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8840;
    wire N__8831;
    wire N__8828;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8824;
    wire N__8823;
    wire N__8812;
    wire N__8809;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8797;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8758;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8707;
    wire N__8704;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8689;
    wire N__8686;
    wire N__8681;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8668;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8650;
    wire N__8649;
    wire N__8648;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8632;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8601;
    wire N__8598;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.un350_ci ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_2_2 ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu0.un88_ci_3_cascade_ ;
    wire \uu0.un55_ci_cascade_ ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.un11_l_count_i ;
    wire uart_RXD;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un284_ci ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire vbuf_tx_data_6;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire vbuf_tx_data_0;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \uu2.r_data_wire_2 ;
    wire vbuf_tx_data_2;
    wire \INVuu2.r_data_reg_2C_net ;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire \uu0.un88_ci_3 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.un66_ci ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un4_l_count_14 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.un4_l_count_18_cascade_ ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un4_l_count_11 ;
    wire \uu0.un4_l_count_16 ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un110_ci ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un165_ci_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_is_det_cascade_ ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.vbuf_raddr.un448_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.un404_ci_0 ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.mem0.N_30_i_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \Lab_UT.dispString.m32_ns_1_cascade_ ;
    wire \Lab_UT.sec1Z0Z_3 ;
    wire \Lab_UT.sec2Z0Z_1 ;
    wire \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ;
    wire \Lab_UT.alarmcharZ0Z_5 ;
    wire \Lab_UT.dispString.m35_ns_1_cascade_ ;
    wire \Lab_UT.dispString.dOut_RNO_0Z0Z_1 ;
    wire \Lab_UT.sec2Z0Z_0 ;
    wire \Lab_UT.alarmcharZ0Z_0 ;
    wire \Lab_UT.dispString.N_46 ;
    wire \Lab_UT.min2Z0Z_1 ;
    wire \Lab_UT.min2Z0Z_2 ;
    wire \Lab_UT.sec1Z0Z_2 ;
    wire \Lab_UT.dicLdAStens_0_cascade_ ;
    wire vbuf_tx_data_rdy;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.un143_ci_0 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \resetGen.reset_count_2_0_4 ;
    wire \Lab_UT.three_2_1_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_2 ;
    wire \Lab_UT.didp.countrce3.q_5_2_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_fastZ0Z_2 ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.didp.did_alarmMatch_6_cascade_ ;
    wire \Lab_UT.min2Z0Z_3 ;
    wire \Lab_UT.min1Z0Z_1 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.didp.regrce1.LdASones_0 ;
    wire \buart.Z_rx.valid_0_cascade_ ;
    wire \buart.Z_rx.idle_0_cascade_ ;
    wire \buart.Z_rx.idle_cascade_ ;
    wire \buart.Z_rx.N_27_0_i_cascade_ ;
    wire bfn_4_14_0_;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.ser_clk_cascade_ ;
    wire \buart.Z_tx.uart_busy_0_0 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.un1_bitcount_c3 ;
    wire \uu2.mem0.w_addr_1 ;
    wire clk;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_ ;
    wire \uu2.mem0.w_data_0_1_3 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_33_0 ;
    wire \uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_ ;
    wire \uu2.mem0.N_409 ;
    wire \uu2.N_34_cascade_ ;
    wire \INVuu2.w_addr_displaying_4C_net ;
    wire \Lab_UT.alarmcharZ0Z_1 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \Lab_UT.dispString.m40_ns_1 ;
    wire \Lab_UT.min1Z0Z_3 ;
    wire \Lab_UT.dispString.N_77_cascade_ ;
    wire \Lab_UT.dispString.N_80 ;
    wire \Lab_UT.sec2Z0Z_3 ;
    wire \Lab_UT.dispString.N_86_cascade_ ;
    wire \Lab_UT.dispString.N_89 ;
    wire \Lab_UT.min2Z0Z_0 ;
    wire \Lab_UT.dispString.m49_ns_1 ;
    wire \Lab_UT.sec1Z0Z_0 ;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire L3_tx_data_5;
    wire L3_tx_data_4;
    wire \Lab_UT.min1Z0Z_0 ;
    wire \Lab_UT.dispString.m25_ns_1 ;
    wire \Lab_UT.min1Z0Z_2 ;
    wire \Lab_UT.dispString.N_65 ;
    wire \Lab_UT.alarmcharZ0Z_6 ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.alarmcharZ0Z_2 ;
    wire \Lab_UT.sec2Z0Z_2 ;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.N_68 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_5 ;
    wire \Lab_UT.didp.did_alarmMatch_11 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ;
    wire \Lab_UT.didp.q_fast_0 ;
    wire \Lab_UT.didp.countrce2.un20_qPone ;
    wire \Lab_UT.didp.countrce2.q_5_3_cascade_ ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.didp.countrce2.q_fastZ0Z_3 ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.didp.countrce2.q_5_3 ;
    wire \Lab_UT.didp.did_alarmMatch_2 ;
    wire \Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_ ;
    wire \Lab_UT.didp.did_alarmMatch_12 ;
    wire \Lab_UT.three_2_0_cascade_ ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.didp.did_alarmMatch_3 ;
    wire \Lab_UT.didp.countrce2.q_fastZ0Z_1 ;
    wire \Lab_UT.didp.countrce3.q_fastZ0Z_1 ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_3_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_fastZ0Z_3 ;
    wire \Lab_UT.didp.q_fast_3 ;
    wire \Lab_UT.didp.countrce3.did_alarmMatch_0 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.dicLdAMones_0_cascade_ ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.dicLdAMones_0 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \resetGen.escKeyZ0Z_5 ;
    wire \resetGen.escKeyZ0Z_4_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.sample ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.startbit_cascade_ ;
    wire bu_rx_data_rdy;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \Lab_UT.didp.countrce2.q_5_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire bfn_6_2_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \uu2.un3_w_addr_user_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.mem0.w_addr_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_44 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_33_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_43 ;
    wire \uu2.N_34 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_42 ;
    wire \uu2.N_49 ;
    wire \uu2.N_57_cascade_ ;
    wire \uu2.w_data_i_a3_0_5 ;
    wire \uu2.mem0.w_data_0_a3_0_6_cascade_ ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.w_data_displaying_2_i_a2_i_a2_0_0 ;
    wire \Lab_UT.alarmcharZ0Z_4 ;
    wire L3_tx_data_6;
    wire L3_tx_data_3;
    wire L3_tx_data_0;
    wire \uu2.un1_w_user_crZ0Z_4 ;
    wire uu2_un1_w_user_cr_0_cascade_;
    wire L3_tx_data_2;
    wire \uu2.mem0.w_data_2 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_ ;
    wire \INVuu2.bitmap_308C_net ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.dictrl.G_64 ;
    wire \Lab_UT.alarmMatch ;
    wire \Lab_UT.dictrl.idle_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ;
    wire \Lab_UT.alarmchar9 ;
    wire \Lab_UT.alarmchar10 ;
    wire \Lab_UT.alarmchar10_i_2 ;
    wire \Lab_UT.dictrl.alarmstateZ0Z_0 ;
    wire \Lab_UT.dictrl.next_alarmstate_1_0 ;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z_0 ;
    wire \Lab_UT.dictrl.next_alarmstate_1_1 ;
    wire \Lab_UT.dictrl.alarmstate_i_3_0 ;
    wire \Lab_UT.dictrl.alarmstateZ0Z_1 ;
    wire \Lab_UT.alarmchar_2_1_1 ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.didp.countrce2.q_5_1 ;
    wire \Lab_UT.didp.countrce2.q_5_2 ;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.didp.countrce3.q_5_1 ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.di_Stens_0 ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.didp.countrce3.q_5_3 ;
    wire \Lab_UT.didp.q_fast_1 ;
    wire \Lab_UT.didp.countrce4.q_5_1 ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.three_2_2_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_5_2_cascade_ ;
    wire \Lab_UT.didp.reset_12_3_3_cascade_ ;
    wire \Lab_UT.didp.reset_12_1_3_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.countrce4.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_5_3 ;
    wire \Lab_UT.didp.countrce4.q_5_0 ;
    wire uu0_sec_clkD;
    wire \Lab_UT.didp.regrce4.LdAMtens_0 ;
    wire \Lab_UT.didp.ce_11_0_2 ;
    wire \Lab_UT.didp.un26_ce_0_cascade_ ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.ce_12_0_3_cascade_ ;
    wire \Lab_UT.didp.un26_ce_0 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.nine_0 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.nine ;
    wire \Lab_UT.five ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_6_13_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \Lab_UT.dictrl.g2_0_1_0_cascade_ ;
    wire bu_rx_data_fast_6;
    wire bu_rx_data_fast_7;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \Lab_UT.dictrl.g2_1_0_0 ;
    wire \INVuu2.w_addr_user_5C_net ;
    wire \uu2.un1_w_user_lf_0_0 ;
    wire \uu2.un1_w_user_lfZ0Z_4 ;
    wire \uu2.un20_w_addr_userZ0Z_1 ;
    wire \uu2.un3_w_addr_user ;
    wire \uu2.un20_w_addr_userZ0Z_1_cascade_ ;
    wire \uu2.w_addr_user_RNI43E87Z0Z_2_cascade_ ;
    wire \uu2.un28_w_addr_user_i ;
    wire \INVuu2.w_addr_user_0C_net ;
    wire \uu2.un3_w_addr_user_5 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.un426_ci_3_cascade_ ;
    wire \uu2.un426_ci_3 ;
    wire \uu2.un404_ci ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.w_addr_user_RNI43E87Z0Z_2 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_42 ;
    wire \INVuu2.w_addr_displaying_nesr_8C_net ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.vbuf_w_addr_user.un448_ci_0 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_0 ;
    wire \INVuu2.bitmap_40C_net ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.bitmap_pmux_sn_N_11_cascade_ ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.N_97_cascade_ ;
    wire \uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2 ;
    wire \Lab_UT.dictrl.next_alarmstate_1 ;
    wire \Lab_UT.dictrl.next_alarmstate_0_0 ;
    wire \Lab_UT.dictrl.un1_next_alarmstate21_0 ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.sec1Z0Z_1 ;
    wire rst;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.escKeyZ0 ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_6 ;
    wire o_One_Sec_Pulse;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \INVuu2.bitmap_93C_net ;
    wire \Lab_UT.bcd2segment3.segment_0Z0Z_0 ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.di_Mones_3 ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \INVuu2.bitmap_296C_net ;
    wire \Lab_UT.didp.countrce1.q_5_0_cascade_ ;
    wire \Lab_UT.three_2 ;
    wire \Lab_UT.didp.countrce1.q_5_2_cascade_ ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.didp.countrce1.q_5_3_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_1 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_ ;
    wire \Lab_UT.LdSones ;
    wire \Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_ ;
    wire \Lab_UT.dicLdSones_1 ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_i_a3_2 ;
    wire \Lab_UT.dictrl.g3_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_a3_2 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.dictrl.g0_1_2_0_cascade_ ;
    wire \Lab_UT.dictrl.N_29_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_30_0 ;
    wire \Lab_UT.dictrl.N_30_0_cascade_ ;
    wire \Lab_UT.dictrl.i6_mux_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.dicLdAMones_0_sx_cascade_ ;
    wire \Lab_UT.dicLdAMones_1 ;
    wire \Lab_UT.dictrl.g0_1_3 ;
    wire \Lab_UT.dictrl.g2_1_0_1_cascade_ ;
    wire \Lab_UT.dictrl.N_7_1_0 ;
    wire bu_rx_data_fast_4;
    wire \Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.next_state18_1_0 ;
    wire \Lab_UT.dictrl.g1_0_1_cascade_ ;
    wire \Lab_UT.dictrl.g2_1 ;
    wire bu_rx_data_fast_5;
    wire bu_rx_data_fast_3;
    wire \uu2.mem0.N_98_0_cascade_ ;
    wire \uu2.mem0.G_11_0_0_a3_0_2 ;
    wire \uu2.mem0.N_62_cascade_ ;
    wire \uu2.mem0.N_36 ;
    wire \uu2.mem0.N_9_cascade_ ;
    wire \uu2.bitmap_pmux_26_bm_1 ;
    wire \uu2.bitmap_RNI31F32Z0Z_34_cascade_ ;
    wire \uu2.w_addr_displaying_RNIBICU6_0Z0Z_2 ;
    wire \uu2.N_401_cascade_ ;
    wire \uu2.w_addr_displaying_RNIBICU6Z0Z_2 ;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.N_99_cascade_ ;
    wire \uu2.bitmap_RNI2Q8F1Z0Z_111 ;
    wire \uu2.bitmap_pmux_sn_N_15 ;
    wire \uu2.bitmap_pmux_sn_N_54_mux ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_fast_nesr_3C_net ;
    wire \uu2.N_31_0 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.N_98_cascade_ ;
    wire \uu2.bitmap_RNI04AD1Z0Z_314 ;
    wire \INVuu2.bitmap_90C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.N_383 ;
    wire L3_tx_data_rdy;
    wire uu2_un1_w_user_cr_0;
    wire \uu2.N_57 ;
    wire \uu2.N_38 ;
    wire \uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \INVuu2.w_addr_displaying_fast_7C_net ;
    wire \Lab_UT.bcd2segment3.segment_0Z0Z_2 ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_4 ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_6 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \Lab_UT.bcd2segment3.segment_0Z0Z_1 ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_5 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \INVuu2.bitmap_203C_net ;
    wire \Lab_UT.LdASones ;
    wire \Lab_UT.LdASones_cascade_ ;
    wire \Lab_UT.LdSones_i_3 ;
    wire \Lab_UT.dicRun_2 ;
    wire \Lab_UT.didp.ce_9_0_0 ;
    wire \Lab_UT.dicRun_2_cascade_ ;
    wire oneSecStrb;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.dictrl.N_11_0 ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_1 ;
    wire \Lab_UT.dictrl.g0_0_i_a3_3_1 ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_3_0 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_4 ;
    wire \Lab_UT.dictrl.N_9_0 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_ ;
    wire bu_rx_data_0;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z4 ;
    wire \Lab_UT.dictrl.N_5_cascade_ ;
    wire \Lab_UT.dictrl.N_10_0 ;
    wire \Lab_UT.dictrl.g0_0_0_o4_0 ;
    wire \Lab_UT.dictrl.N_3_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_a3_2_0 ;
    wire \Lab_UT.dictrl.g0_0_i_o4_0 ;
    wire \Lab_UT.dictrl.g0_1Z0Z_2 ;
    wire \Lab_UT.dictrl.next_state18_0 ;
    wire \Lab_UT.dictrl.next_state18_0_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_7_0 ;
    wire \Lab_UT.dictrl.N_11 ;
    wire \Lab_UT.dictrl.g2_2_0 ;
    wire \Lab_UT.dictrl.next_alarmstate4Z0Z_3 ;
    wire \Lab_UT.dictrl.next_alarmstate4Z0Z_0 ;
    wire \Lab_UT.dictrl.g2_1_2 ;
    wire \Lab_UT.dictrl.g1_5_1_cascade_ ;
    wire \Lab_UT.dictrl.g2_3 ;
    wire \Lab_UT.dictrl.g0Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_3_cascade_ ;
    wire bu_rx_data_5_rep1;
    wire \Lab_UT.dictrl.next_state12_0 ;
    wire bu_rx_data_6_rep1;
    wire \Lab_UT.dictrl.g0_8Z0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.g2_1_3 ;
    wire bu_rx_data_1_rep1;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_28 ;
    wire \uu2.mem0.N_44 ;
    wire \uu2.mem0.N_41_cascade_ ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.bitmap_pmux_sn_N_36 ;
    wire \uu2.mem0.N_24_i_cascade_ ;
    wire \uu2.N_406 ;
    wire \uu2.mem0.N_45 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.mem0.G_11_0_0_a2_3_4 ;
    wire N_272_mux;
    wire \uu2.mem0.G_11_0_0_a2_3_5_cascade_ ;
    wire L3_tx_data_1;
    wire \uu2.mem0.G_11_0_0_0 ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_1 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_5 ;
    wire \Lab_UT.bcd2segment2.segmentUQ_0_4 ;
    wire \Lab_UT.bcd2segment2.segment_0Z0Z_2 ;
    wire \INVuu2.bitmap_87C_net ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmap_pmux_17_ns_1_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.N_104_cascade_ ;
    wire \uu2.mem0.G_11_0_0_a3_5_0_cascade_ ;
    wire \uu2.mem0.N_40 ;
    wire \uu2.mem0.N_30 ;
    wire \uu2.w_addr_displaying_2_repZ0Z1 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_41 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.w_addr_displaying_RNIVAPV6Z0Z_5 ;
    wire \INVuu2.w_addr_displaying_2_rep1C_net ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.bitmap_pmux_20_ns_1_cascade_ ;
    wire \uu2.mem0.N_108 ;
    wire \INVuu2.bitmap_194C_net ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.bitmap_pmux_20_ns_1 ;
    wire \uu2.mem0.N_108_0_cascade_ ;
    wire \uu2.mem0.N_404_0 ;
    wire \uu2.mem0.bitmap_pmux_16_ns_1_cascade_ ;
    wire \uu2.N_30_i ;
    wire \uu2.mem0.N_22_cascade_ ;
    wire \uu2.mem0.G_11_0_0_a3_6_0 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_ ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.N_30_i_1 ;
    wire \uu2.mem0.N_22_0_cascade_ ;
    wire \uu2.N_104 ;
    wire \uu2.mem0.bitmap_pmux_27_ns_1_0 ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.mem0.N_109 ;
    wire \uu2.bitmap_pmux_19_ns_1 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.mem0.N_109_0 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_3 ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_2 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_5 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_6 ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_0 ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_1 ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \INVuu2.bitmap_218C_net ;
    wire \Lab_UT.dictrl.N_14_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_i_a3_0_3 ;
    wire \Lab_UT.dictrl.N_7_cascade_ ;
    wire \Lab_UT.dictrl.N_13_0_cascade_ ;
    wire \Lab_UT.dictrl.N_6_cascade_ ;
    wire \Lab_UT.LdStens ;
    wire \Lab_UT.state_i_3_2 ;
    wire \Lab_UT.LdStens_i_3 ;
    wire \Lab_UT.didp.ce_10_0_1 ;
    wire \Lab_UT.dictrl.m27_1 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_0 ;
    wire \Lab_UT.dictrl.N_19_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.N_19 ;
    wire \Lab_UT.dictrl.N_11_0_0 ;
    wire \Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_5_RNOZ0Z_1 ;
    wire \Lab_UT.dicRun_1 ;
    wire \Lab_UT.dictrl.N_10 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_2 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_ ;
    wire \Lab_UT.dictrl.N_5 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_3 ;
    wire \Lab_UT.dictrl.i6_mux ;
    wire \Lab_UT.dictrl.N_15_0_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1 ;
    wire \Lab_UT.dictrl.state_i_3Z0Z_0 ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.dictrl.g0_6_o3_2_0_cascade_ ;
    wire \Lab_UT.dictrl.N_5_0_cascade_ ;
    wire \Lab_UT.dictrl.g1_3_0 ;
    wire \Lab_UT.dictrl.g2_2 ;
    wire \Lab_UT.dictrl.N_16_0_0 ;
    wire \Lab_UT.dictrl.g0_i_a3_0_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a3_0_6_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a3_0_5 ;
    wire \Lab_UT.dictrl.N_3 ;
    wire \Lab_UT.dictrl.g1_4 ;
    wire \Lab_UT.dictrl.gZ0Z1 ;
    wire \Lab_UT.dictrl.next_state12_1 ;
    wire \Lab_UT.dictrl.next_state32Z0Z_4 ;
    wire \Lab_UT.dictrl.g1Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.N_13_0_0 ;
    wire \Lab_UT.dictrl.g1_2_2_cascade_ ;
    wire \Lab_UT.dictrl.g2_1_1 ;
    wire \Lab_UT.dictrl.g2_0 ;
    wire \Lab_UT.dictrl.g1_2_3 ;
    wire \Lab_UT.dictrl.g0_1Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_i_a3_4 ;
    wire bu_rx_data_4_rep1;
    wire bu_rx_data_7_rep1;
    wire \Lab_UT.dictrl.g1_4_0 ;
    wire bu_rx_data_2_rep1;
    wire bu_rx_data_fast_2;
    wire bu_rx_data_3;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_2;
    wire bu_rx_data_3_rep1;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \INVuu2.bitmap_34C_net ;
    wire \Lab_UT.bcd2segment4.segment_0Z0Z_2 ;
    wire \Lab_UT.bcd2segment4.segmentUQ_0_4 ;
    wire \Lab_UT.bcd2segment4.segmentUQ_0_5 ;
    wire \Lab_UT.bcd2segment4.segmentUQ_0_6 ;
    wire \Lab_UT.bcd2segment4.segment_0Z0Z_0 ;
    wire \Lab_UT.bcd2segment4.segment_0Z0Z_1 ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_ ;
    wire \Lab_UT.Run ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \Lab_UT.dictrl.N_39_mux ;
    wire \Lab_UT.dictrl.g0_0_a3_2 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_1 ;
    wire \Lab_UT.dictrl.un1_next_state66_0 ;
    wire \Lab_UT.dictrl.g0_0_i_a3_1 ;
    wire \Lab_UT.dicLdAStens_0 ;
    wire \Lab_UT.dictrl.N_40_mux ;
    wire \Lab_UT.state_3 ;
    wire \Lab_UT.dictrl.N_13_cascade_ ;
    wire \Lab_UT.dictrl.N_16 ;
    wire \Lab_UT.dictrl.state_fast_3 ;
    wire bu_rx_data_2_rep2;
    wire \Lab_UT.dictrl.N_15 ;
    wire \Lab_UT.dictrl.next_state12 ;
    wire \Lab_UT.dictrl.stateZ0Z_2 ;
    wire \Lab_UT.dictrl.N_21_cascade_ ;
    wire \Lab_UT.dictrl.next_state_latmux_0_1 ;
    wire \Lab_UT.dictrl.next_state18 ;
    wire bu_rx_data_1_rep2;
    wire \Lab_UT.dictrl.g1_5_0 ;
    wire \Lab_UT.state_1 ;
    wire \Lab_UT.dictrl.N_23 ;
    wire \Lab_UT.dictrl.N_30 ;
    wire \Lab_UT.dictrl.next_state5_3_cascade_ ;
    wire \Lab_UT.dictrl.next_state32Z0Z_1 ;
    wire \Lab_UT.dictrl.N_18 ;
    wire \Lab_UT.dictrl.state_3_rep1 ;
    wire \Lab_UT.dictrl.m17_1 ;
    wire \Lab_UT.state_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z32 ;
    wire \Lab_UT.dictrl.N_29_0 ;
    wire bu_rx_data_fast_0;
    wire \Lab_UT.dictrl.g1_5_cascade_ ;
    wire \Lab_UT.dictrl.g1_6 ;
    wire \Lab_UT.dictrl.g1_0_0 ;
    wire \Lab_UT.dictrl.state_3_rep2 ;
    wire \Lab_UT.dictrl.g0_i_a3_3 ;
    wire bu_rx_data_7;
    wire bu_rx_data_3_rep2;
    wire bu_rx_data_6;
    wire bu_rx_data_1;
    wire bu_rx_data_0_rep1;
    wire bu_rx_data_5;
    wire bu_rx_data_4;
    wire _gnd_net_;
    wire clk_g;
    wire \buart.Z_rx.sample_g ;
    wire rst_g;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__8588),
            .RESETB(N__12671),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__10175,N__10151,N__10046,N__10079,N__10112,N__9923,N__10022,N__9989,N__9959}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__12251,N__14003,N__14021,N__11153,N__10931,N__11207,N__12398,N__10985,N__12236}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__12542,dangling_wire_31,N__10226,dangling_wire_32,N__10238,dangling_wire_33,N__10217,dangling_wire_34,N__12416,dangling_wire_35,N__16823,dangling_wire_36,N__10232}),
            .RCLKE(),
            .RCLK(N__22354),
            .RE(N__12664),
            .WCLKE(N__10952),
            .WCLK(N__22353),
            .WE(N__10948));
    IO_PAD led_obuft_3_iopad (
            .OE(N__23331),
            .DIN(N__23330),
            .DOUT(N__23329),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__23331),
            .PADOUT(N__23330),
            .PADIN(N__23329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__23322),
            .DIN(N__23321),
            .DOUT(N__23320),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__23322),
            .PADOUT(N__23321),
            .PADIN(N__23320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__23313),
            .DIN(N__23312),
            .DOUT(N__23311),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__23313),
            .PADOUT(N__23312),
            .PADIN(N__23311),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__22321),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__23304),
            .DIN(N__23303),
            .DOUT(N__23302),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__23304),
            .PADOUT(N__23303),
            .PADIN(N__23302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__23295),
            .DIN(N__23294),
            .DOUT(N__23293),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__23295),
            .PADOUT(N__23294),
            .PADIN(N__23293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__23286),
            .DIN(N__23285),
            .DOUT(N__23284),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__23286),
            .PADOUT(N__23285),
            .PADIN(N__23284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__23277),
            .DIN(N__23276),
            .DOUT(N__23275),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__23277),
            .PADOUT(N__23276),
            .PADIN(N__23275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__23268),
            .DIN(N__23267),
            .DOUT(N__23266),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__23268),
            .PADOUT(N__23267),
            .PADIN(N__23266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9314),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__23259),
            .DIN(N__23258),
            .DOUT(N__23257),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__23259),
            .PADOUT(N__23258),
            .PADIN(N__23257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__23250),
            .DIN(N__23249),
            .DOUT(N__23248),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__23250),
            .PADOUT(N__23249),
            .PADIN(N__23248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__5612 (
            .O(N__23231),
            .I(\Lab_UT.dictrl.g1_5_cascade_ ));
    InMux I__5611 (
            .O(N__23228),
            .I(N__23225));
    LocalMux I__5610 (
            .O(N__23225),
            .I(\Lab_UT.dictrl.g1_6 ));
    InMux I__5609 (
            .O(N__23222),
            .I(N__23219));
    LocalMux I__5608 (
            .O(N__23219),
            .I(N__23216));
    Span4Mux_h I__5607 (
            .O(N__23216),
            .I(N__23213));
    Odrv4 I__5606 (
            .O(N__23213),
            .I(\Lab_UT.dictrl.g1_0_0 ));
    InMux I__5605 (
            .O(N__23210),
            .I(N__23206));
    InMux I__5604 (
            .O(N__23209),
            .I(N__23199));
    LocalMux I__5603 (
            .O(N__23206),
            .I(N__23189));
    InMux I__5602 (
            .O(N__23205),
            .I(N__23182));
    InMux I__5601 (
            .O(N__23204),
            .I(N__23182));
    InMux I__5600 (
            .O(N__23203),
            .I(N__23182));
    InMux I__5599 (
            .O(N__23202),
            .I(N__23178));
    LocalMux I__5598 (
            .O(N__23199),
            .I(N__23175));
    CascadeMux I__5597 (
            .O(N__23198),
            .I(N__23171));
    CascadeMux I__5596 (
            .O(N__23197),
            .I(N__23167));
    InMux I__5595 (
            .O(N__23196),
            .I(N__23160));
    InMux I__5594 (
            .O(N__23195),
            .I(N__23160));
    InMux I__5593 (
            .O(N__23194),
            .I(N__23160));
    InMux I__5592 (
            .O(N__23193),
            .I(N__23155));
    InMux I__5591 (
            .O(N__23192),
            .I(N__23155));
    Span4Mux_h I__5590 (
            .O(N__23189),
            .I(N__23150));
    LocalMux I__5589 (
            .O(N__23182),
            .I(N__23150));
    InMux I__5588 (
            .O(N__23181),
            .I(N__23147));
    LocalMux I__5587 (
            .O(N__23178),
            .I(N__23144));
    Span4Mux_v I__5586 (
            .O(N__23175),
            .I(N__23141));
    InMux I__5585 (
            .O(N__23174),
            .I(N__23138));
    InMux I__5584 (
            .O(N__23171),
            .I(N__23135));
    InMux I__5583 (
            .O(N__23170),
            .I(N__23130));
    InMux I__5582 (
            .O(N__23167),
            .I(N__23130));
    LocalMux I__5581 (
            .O(N__23160),
            .I(N__23125));
    LocalMux I__5580 (
            .O(N__23155),
            .I(N__23125));
    Span4Mux_h I__5579 (
            .O(N__23150),
            .I(N__23122));
    LocalMux I__5578 (
            .O(N__23147),
            .I(N__23117));
    Span4Mux_h I__5577 (
            .O(N__23144),
            .I(N__23117));
    Span4Mux_h I__5576 (
            .O(N__23141),
            .I(N__23108));
    LocalMux I__5575 (
            .O(N__23138),
            .I(N__23108));
    LocalMux I__5574 (
            .O(N__23135),
            .I(N__23108));
    LocalMux I__5573 (
            .O(N__23130),
            .I(N__23108));
    Span12Mux_s10_h I__5572 (
            .O(N__23125),
            .I(N__23105));
    Odrv4 I__5571 (
            .O(N__23122),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv4 I__5570 (
            .O(N__23117),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv4 I__5569 (
            .O(N__23108),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv12 I__5568 (
            .O(N__23105),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    InMux I__5567 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__5566 (
            .O(N__23093),
            .I(N__23090));
    Odrv4 I__5565 (
            .O(N__23090),
            .I(\Lab_UT.dictrl.g0_i_a3_3 ));
    CascadeMux I__5564 (
            .O(N__23087),
            .I(N__23080));
    CascadeMux I__5563 (
            .O(N__23086),
            .I(N__23074));
    InMux I__5562 (
            .O(N__23085),
            .I(N__23069));
    InMux I__5561 (
            .O(N__23084),
            .I(N__23066));
    InMux I__5560 (
            .O(N__23083),
            .I(N__23061));
    InMux I__5559 (
            .O(N__23080),
            .I(N__23061));
    InMux I__5558 (
            .O(N__23079),
            .I(N__23058));
    InMux I__5557 (
            .O(N__23078),
            .I(N__23055));
    InMux I__5556 (
            .O(N__23077),
            .I(N__23052));
    InMux I__5555 (
            .O(N__23074),
            .I(N__23047));
    InMux I__5554 (
            .O(N__23073),
            .I(N__23047));
    InMux I__5553 (
            .O(N__23072),
            .I(N__23042));
    LocalMux I__5552 (
            .O(N__23069),
            .I(N__23035));
    LocalMux I__5551 (
            .O(N__23066),
            .I(N__23035));
    LocalMux I__5550 (
            .O(N__23061),
            .I(N__23035));
    LocalMux I__5549 (
            .O(N__23058),
            .I(N__23030));
    LocalMux I__5548 (
            .O(N__23055),
            .I(N__23025));
    LocalMux I__5547 (
            .O(N__23052),
            .I(N__23025));
    LocalMux I__5546 (
            .O(N__23047),
            .I(N__23022));
    InMux I__5545 (
            .O(N__23046),
            .I(N__23017));
    InMux I__5544 (
            .O(N__23045),
            .I(N__23017));
    LocalMux I__5543 (
            .O(N__23042),
            .I(N__23014));
    Span4Mux_v I__5542 (
            .O(N__23035),
            .I(N__23011));
    InMux I__5541 (
            .O(N__23034),
            .I(N__23008));
    InMux I__5540 (
            .O(N__23033),
            .I(N__23005));
    Span4Mux_v I__5539 (
            .O(N__23030),
            .I(N__23002));
    Span4Mux_h I__5538 (
            .O(N__23025),
            .I(N__22999));
    Span4Mux_v I__5537 (
            .O(N__23022),
            .I(N__22994));
    LocalMux I__5536 (
            .O(N__23017),
            .I(N__22994));
    Span4Mux_s2_v I__5535 (
            .O(N__23014),
            .I(N__22989));
    Span4Mux_h I__5534 (
            .O(N__23011),
            .I(N__22989));
    LocalMux I__5533 (
            .O(N__23008),
            .I(bu_rx_data_7));
    LocalMux I__5532 (
            .O(N__23005),
            .I(bu_rx_data_7));
    Odrv4 I__5531 (
            .O(N__23002),
            .I(bu_rx_data_7));
    Odrv4 I__5530 (
            .O(N__22999),
            .I(bu_rx_data_7));
    Odrv4 I__5529 (
            .O(N__22994),
            .I(bu_rx_data_7));
    Odrv4 I__5528 (
            .O(N__22989),
            .I(bu_rx_data_7));
    InMux I__5527 (
            .O(N__22976),
            .I(N__22966));
    CascadeMux I__5526 (
            .O(N__22975),
            .I(N__22962));
    InMux I__5525 (
            .O(N__22974),
            .I(N__22956));
    InMux I__5524 (
            .O(N__22973),
            .I(N__22953));
    CascadeMux I__5523 (
            .O(N__22972),
            .I(N__22949));
    CascadeMux I__5522 (
            .O(N__22971),
            .I(N__22946));
    InMux I__5521 (
            .O(N__22970),
            .I(N__22941));
    InMux I__5520 (
            .O(N__22969),
            .I(N__22941));
    LocalMux I__5519 (
            .O(N__22966),
            .I(N__22938));
    InMux I__5518 (
            .O(N__22965),
            .I(N__22933));
    InMux I__5517 (
            .O(N__22962),
            .I(N__22933));
    InMux I__5516 (
            .O(N__22961),
            .I(N__22930));
    InMux I__5515 (
            .O(N__22960),
            .I(N__22925));
    InMux I__5514 (
            .O(N__22959),
            .I(N__22925));
    LocalMux I__5513 (
            .O(N__22956),
            .I(N__22920));
    LocalMux I__5512 (
            .O(N__22953),
            .I(N__22920));
    InMux I__5511 (
            .O(N__22952),
            .I(N__22917));
    InMux I__5510 (
            .O(N__22949),
            .I(N__22914));
    InMux I__5509 (
            .O(N__22946),
            .I(N__22911));
    LocalMux I__5508 (
            .O(N__22941),
            .I(N__22904));
    Span4Mux_h I__5507 (
            .O(N__22938),
            .I(N__22904));
    LocalMux I__5506 (
            .O(N__22933),
            .I(N__22904));
    LocalMux I__5505 (
            .O(N__22930),
            .I(N__22901));
    LocalMux I__5504 (
            .O(N__22925),
            .I(N__22898));
    Span4Mux_h I__5503 (
            .O(N__22920),
            .I(N__22895));
    LocalMux I__5502 (
            .O(N__22917),
            .I(N__22886));
    LocalMux I__5501 (
            .O(N__22914),
            .I(N__22886));
    LocalMux I__5500 (
            .O(N__22911),
            .I(N__22886));
    Span4Mux_v I__5499 (
            .O(N__22904),
            .I(N__22886));
    Odrv4 I__5498 (
            .O(N__22901),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5497 (
            .O(N__22898),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5496 (
            .O(N__22895),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5495 (
            .O(N__22886),
            .I(bu_rx_data_3_rep2));
    InMux I__5494 (
            .O(N__22877),
            .I(N__22872));
    InMux I__5493 (
            .O(N__22876),
            .I(N__22866));
    CascadeMux I__5492 (
            .O(N__22875),
            .I(N__22859));
    LocalMux I__5491 (
            .O(N__22872),
            .I(N__22856));
    CascadeMux I__5490 (
            .O(N__22871),
            .I(N__22853));
    InMux I__5489 (
            .O(N__22870),
            .I(N__22848));
    InMux I__5488 (
            .O(N__22869),
            .I(N__22848));
    LocalMux I__5487 (
            .O(N__22866),
            .I(N__22845));
    InMux I__5486 (
            .O(N__22865),
            .I(N__22842));
    InMux I__5485 (
            .O(N__22864),
            .I(N__22839));
    InMux I__5484 (
            .O(N__22863),
            .I(N__22834));
    InMux I__5483 (
            .O(N__22862),
            .I(N__22834));
    InMux I__5482 (
            .O(N__22859),
            .I(N__22831));
    Span4Mux_s2_h I__5481 (
            .O(N__22856),
            .I(N__22828));
    InMux I__5480 (
            .O(N__22853),
            .I(N__22821));
    LocalMux I__5479 (
            .O(N__22848),
            .I(N__22814));
    Span4Mux_h I__5478 (
            .O(N__22845),
            .I(N__22814));
    LocalMux I__5477 (
            .O(N__22842),
            .I(N__22814));
    LocalMux I__5476 (
            .O(N__22839),
            .I(N__22809));
    LocalMux I__5475 (
            .O(N__22834),
            .I(N__22809));
    LocalMux I__5474 (
            .O(N__22831),
            .I(N__22804));
    Span4Mux_h I__5473 (
            .O(N__22828),
            .I(N__22804));
    InMux I__5472 (
            .O(N__22827),
            .I(N__22801));
    InMux I__5471 (
            .O(N__22826),
            .I(N__22798));
    InMux I__5470 (
            .O(N__22825),
            .I(N__22793));
    InMux I__5469 (
            .O(N__22824),
            .I(N__22793));
    LocalMux I__5468 (
            .O(N__22821),
            .I(N__22788));
    Span4Mux_h I__5467 (
            .O(N__22814),
            .I(N__22788));
    Span4Mux_v I__5466 (
            .O(N__22809),
            .I(N__22785));
    Span4Mux_h I__5465 (
            .O(N__22804),
            .I(N__22782));
    LocalMux I__5464 (
            .O(N__22801),
            .I(bu_rx_data_6));
    LocalMux I__5463 (
            .O(N__22798),
            .I(bu_rx_data_6));
    LocalMux I__5462 (
            .O(N__22793),
            .I(bu_rx_data_6));
    Odrv4 I__5461 (
            .O(N__22788),
            .I(bu_rx_data_6));
    Odrv4 I__5460 (
            .O(N__22785),
            .I(bu_rx_data_6));
    Odrv4 I__5459 (
            .O(N__22782),
            .I(bu_rx_data_6));
    InMux I__5458 (
            .O(N__22769),
            .I(N__22761));
    InMux I__5457 (
            .O(N__22768),
            .I(N__22756));
    InMux I__5456 (
            .O(N__22767),
            .I(N__22752));
    InMux I__5455 (
            .O(N__22766),
            .I(N__22749));
    InMux I__5454 (
            .O(N__22765),
            .I(N__22744));
    InMux I__5453 (
            .O(N__22764),
            .I(N__22738));
    LocalMux I__5452 (
            .O(N__22761),
            .I(N__22733));
    InMux I__5451 (
            .O(N__22760),
            .I(N__22728));
    InMux I__5450 (
            .O(N__22759),
            .I(N__22728));
    LocalMux I__5449 (
            .O(N__22756),
            .I(N__22724));
    InMux I__5448 (
            .O(N__22755),
            .I(N__22721));
    LocalMux I__5447 (
            .O(N__22752),
            .I(N__22716));
    LocalMux I__5446 (
            .O(N__22749),
            .I(N__22716));
    InMux I__5445 (
            .O(N__22748),
            .I(N__22713));
    InMux I__5444 (
            .O(N__22747),
            .I(N__22710));
    LocalMux I__5443 (
            .O(N__22744),
            .I(N__22707));
    InMux I__5442 (
            .O(N__22743),
            .I(N__22702));
    InMux I__5441 (
            .O(N__22742),
            .I(N__22697));
    InMux I__5440 (
            .O(N__22741),
            .I(N__22697));
    LocalMux I__5439 (
            .O(N__22738),
            .I(N__22694));
    InMux I__5438 (
            .O(N__22737),
            .I(N__22691));
    InMux I__5437 (
            .O(N__22736),
            .I(N__22688));
    Span4Mux_s3_v I__5436 (
            .O(N__22733),
            .I(N__22685));
    LocalMux I__5435 (
            .O(N__22728),
            .I(N__22682));
    InMux I__5434 (
            .O(N__22727),
            .I(N__22679));
    Span4Mux_v I__5433 (
            .O(N__22724),
            .I(N__22672));
    LocalMux I__5432 (
            .O(N__22721),
            .I(N__22672));
    Span4Mux_v I__5431 (
            .O(N__22716),
            .I(N__22672));
    LocalMux I__5430 (
            .O(N__22713),
            .I(N__22665));
    LocalMux I__5429 (
            .O(N__22710),
            .I(N__22665));
    Span4Mux_v I__5428 (
            .O(N__22707),
            .I(N__22665));
    InMux I__5427 (
            .O(N__22706),
            .I(N__22660));
    InMux I__5426 (
            .O(N__22705),
            .I(N__22660));
    LocalMux I__5425 (
            .O(N__22702),
            .I(N__22655));
    LocalMux I__5424 (
            .O(N__22697),
            .I(N__22655));
    Span4Mux_s2_h I__5423 (
            .O(N__22694),
            .I(N__22652));
    LocalMux I__5422 (
            .O(N__22691),
            .I(N__22647));
    LocalMux I__5421 (
            .O(N__22688),
            .I(N__22647));
    Span4Mux_h I__5420 (
            .O(N__22685),
            .I(N__22642));
    Span4Mux_v I__5419 (
            .O(N__22682),
            .I(N__22642));
    LocalMux I__5418 (
            .O(N__22679),
            .I(N__22635));
    Span4Mux_v I__5417 (
            .O(N__22672),
            .I(N__22635));
    Span4Mux_v I__5416 (
            .O(N__22665),
            .I(N__22635));
    LocalMux I__5415 (
            .O(N__22660),
            .I(N__22630));
    Span4Mux_h I__5414 (
            .O(N__22655),
            .I(N__22630));
    Span4Mux_h I__5413 (
            .O(N__22652),
            .I(N__22627));
    Odrv12 I__5412 (
            .O(N__22647),
            .I(bu_rx_data_1));
    Odrv4 I__5411 (
            .O(N__22642),
            .I(bu_rx_data_1));
    Odrv4 I__5410 (
            .O(N__22635),
            .I(bu_rx_data_1));
    Odrv4 I__5409 (
            .O(N__22630),
            .I(bu_rx_data_1));
    Odrv4 I__5408 (
            .O(N__22627),
            .I(bu_rx_data_1));
    CascadeMux I__5407 (
            .O(N__22616),
            .I(N__22612));
    CascadeMux I__5406 (
            .O(N__22615),
            .I(N__22606));
    InMux I__5405 (
            .O(N__22612),
            .I(N__22603));
    CascadeMux I__5404 (
            .O(N__22611),
            .I(N__22600));
    InMux I__5403 (
            .O(N__22610),
            .I(N__22592));
    InMux I__5402 (
            .O(N__22609),
            .I(N__22592));
    InMux I__5401 (
            .O(N__22606),
            .I(N__22592));
    LocalMux I__5400 (
            .O(N__22603),
            .I(N__22589));
    InMux I__5399 (
            .O(N__22600),
            .I(N__22586));
    InMux I__5398 (
            .O(N__22599),
            .I(N__22583));
    LocalMux I__5397 (
            .O(N__22592),
            .I(N__22580));
    Span4Mux_h I__5396 (
            .O(N__22589),
            .I(N__22577));
    LocalMux I__5395 (
            .O(N__22586),
            .I(N__22574));
    LocalMux I__5394 (
            .O(N__22583),
            .I(N__22571));
    Span4Mux_h I__5393 (
            .O(N__22580),
            .I(N__22568));
    Odrv4 I__5392 (
            .O(N__22577),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__5391 (
            .O(N__22574),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__5390 (
            .O(N__22571),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__5389 (
            .O(N__22568),
            .I(bu_rx_data_0_rep1));
    InMux I__5388 (
            .O(N__22559),
            .I(N__22553));
    InMux I__5387 (
            .O(N__22558),
            .I(N__22550));
    CascadeMux I__5386 (
            .O(N__22557),
            .I(N__22547));
    InMux I__5385 (
            .O(N__22556),
            .I(N__22541));
    LocalMux I__5384 (
            .O(N__22553),
            .I(N__22536));
    LocalMux I__5383 (
            .O(N__22550),
            .I(N__22536));
    InMux I__5382 (
            .O(N__22547),
            .I(N__22533));
    InMux I__5381 (
            .O(N__22546),
            .I(N__22528));
    InMux I__5380 (
            .O(N__22545),
            .I(N__22524));
    InMux I__5379 (
            .O(N__22544),
            .I(N__22521));
    LocalMux I__5378 (
            .O(N__22541),
            .I(N__22513));
    Span4Mux_v I__5377 (
            .O(N__22536),
            .I(N__22513));
    LocalMux I__5376 (
            .O(N__22533),
            .I(N__22513));
    InMux I__5375 (
            .O(N__22532),
            .I(N__22508));
    InMux I__5374 (
            .O(N__22531),
            .I(N__22508));
    LocalMux I__5373 (
            .O(N__22528),
            .I(N__22505));
    InMux I__5372 (
            .O(N__22527),
            .I(N__22499));
    LocalMux I__5371 (
            .O(N__22524),
            .I(N__22494));
    LocalMux I__5370 (
            .O(N__22521),
            .I(N__22494));
    InMux I__5369 (
            .O(N__22520),
            .I(N__22491));
    Span4Mux_h I__5368 (
            .O(N__22513),
            .I(N__22488));
    LocalMux I__5367 (
            .O(N__22508),
            .I(N__22483));
    Span12Mux_v I__5366 (
            .O(N__22505),
            .I(N__22483));
    InMux I__5365 (
            .O(N__22504),
            .I(N__22476));
    InMux I__5364 (
            .O(N__22503),
            .I(N__22476));
    InMux I__5363 (
            .O(N__22502),
            .I(N__22476));
    LocalMux I__5362 (
            .O(N__22499),
            .I(N__22471));
    Span4Mux_s3_v I__5361 (
            .O(N__22494),
            .I(N__22471));
    LocalMux I__5360 (
            .O(N__22491),
            .I(bu_rx_data_5));
    Odrv4 I__5359 (
            .O(N__22488),
            .I(bu_rx_data_5));
    Odrv12 I__5358 (
            .O(N__22483),
            .I(bu_rx_data_5));
    LocalMux I__5357 (
            .O(N__22476),
            .I(bu_rx_data_5));
    Odrv4 I__5356 (
            .O(N__22471),
            .I(bu_rx_data_5));
    InMux I__5355 (
            .O(N__22460),
            .I(N__22452));
    InMux I__5354 (
            .O(N__22459),
            .I(N__22446));
    InMux I__5353 (
            .O(N__22458),
            .I(N__22443));
    InMux I__5352 (
            .O(N__22457),
            .I(N__22440));
    InMux I__5351 (
            .O(N__22456),
            .I(N__22437));
    InMux I__5350 (
            .O(N__22455),
            .I(N__22431));
    LocalMux I__5349 (
            .O(N__22452),
            .I(N__22427));
    InMux I__5348 (
            .O(N__22451),
            .I(N__22420));
    InMux I__5347 (
            .O(N__22450),
            .I(N__22420));
    InMux I__5346 (
            .O(N__22449),
            .I(N__22420));
    LocalMux I__5345 (
            .O(N__22446),
            .I(N__22416));
    LocalMux I__5344 (
            .O(N__22443),
            .I(N__22409));
    LocalMux I__5343 (
            .O(N__22440),
            .I(N__22409));
    LocalMux I__5342 (
            .O(N__22437),
            .I(N__22409));
    InMux I__5341 (
            .O(N__22436),
            .I(N__22402));
    InMux I__5340 (
            .O(N__22435),
            .I(N__22402));
    InMux I__5339 (
            .O(N__22434),
            .I(N__22402));
    LocalMux I__5338 (
            .O(N__22431),
            .I(N__22399));
    InMux I__5337 (
            .O(N__22430),
            .I(N__22396));
    Span4Mux_h I__5336 (
            .O(N__22427),
            .I(N__22391));
    LocalMux I__5335 (
            .O(N__22420),
            .I(N__22391));
    InMux I__5334 (
            .O(N__22419),
            .I(N__22388));
    Span4Mux_h I__5333 (
            .O(N__22416),
            .I(N__22385));
    Span4Mux_h I__5332 (
            .O(N__22409),
            .I(N__22380));
    LocalMux I__5331 (
            .O(N__22402),
            .I(N__22380));
    Span4Mux_v I__5330 (
            .O(N__22399),
            .I(N__22375));
    LocalMux I__5329 (
            .O(N__22396),
            .I(N__22375));
    Span4Mux_h I__5328 (
            .O(N__22391),
            .I(N__22372));
    LocalMux I__5327 (
            .O(N__22388),
            .I(bu_rx_data_4));
    Odrv4 I__5326 (
            .O(N__22385),
            .I(bu_rx_data_4));
    Odrv4 I__5325 (
            .O(N__22380),
            .I(bu_rx_data_4));
    Odrv4 I__5324 (
            .O(N__22375),
            .I(bu_rx_data_4));
    Odrv4 I__5323 (
            .O(N__22372),
            .I(bu_rx_data_4));
    ClkMux I__5322 (
            .O(N__22361),
            .I(N__22082));
    ClkMux I__5321 (
            .O(N__22360),
            .I(N__22082));
    ClkMux I__5320 (
            .O(N__22359),
            .I(N__22082));
    ClkMux I__5319 (
            .O(N__22358),
            .I(N__22082));
    ClkMux I__5318 (
            .O(N__22357),
            .I(N__22082));
    ClkMux I__5317 (
            .O(N__22356),
            .I(N__22082));
    ClkMux I__5316 (
            .O(N__22355),
            .I(N__22082));
    ClkMux I__5315 (
            .O(N__22354),
            .I(N__22082));
    ClkMux I__5314 (
            .O(N__22353),
            .I(N__22082));
    ClkMux I__5313 (
            .O(N__22352),
            .I(N__22082));
    ClkMux I__5312 (
            .O(N__22351),
            .I(N__22082));
    ClkMux I__5311 (
            .O(N__22350),
            .I(N__22082));
    ClkMux I__5310 (
            .O(N__22349),
            .I(N__22082));
    ClkMux I__5309 (
            .O(N__22348),
            .I(N__22082));
    ClkMux I__5308 (
            .O(N__22347),
            .I(N__22082));
    ClkMux I__5307 (
            .O(N__22346),
            .I(N__22082));
    ClkMux I__5306 (
            .O(N__22345),
            .I(N__22082));
    ClkMux I__5305 (
            .O(N__22344),
            .I(N__22082));
    ClkMux I__5304 (
            .O(N__22343),
            .I(N__22082));
    ClkMux I__5303 (
            .O(N__22342),
            .I(N__22082));
    ClkMux I__5302 (
            .O(N__22341),
            .I(N__22082));
    ClkMux I__5301 (
            .O(N__22340),
            .I(N__22082));
    ClkMux I__5300 (
            .O(N__22339),
            .I(N__22082));
    ClkMux I__5299 (
            .O(N__22338),
            .I(N__22082));
    ClkMux I__5298 (
            .O(N__22337),
            .I(N__22082));
    ClkMux I__5297 (
            .O(N__22336),
            .I(N__22082));
    ClkMux I__5296 (
            .O(N__22335),
            .I(N__22082));
    ClkMux I__5295 (
            .O(N__22334),
            .I(N__22082));
    ClkMux I__5294 (
            .O(N__22333),
            .I(N__22082));
    ClkMux I__5293 (
            .O(N__22332),
            .I(N__22082));
    ClkMux I__5292 (
            .O(N__22331),
            .I(N__22082));
    ClkMux I__5291 (
            .O(N__22330),
            .I(N__22082));
    ClkMux I__5290 (
            .O(N__22329),
            .I(N__22082));
    ClkMux I__5289 (
            .O(N__22328),
            .I(N__22082));
    ClkMux I__5288 (
            .O(N__22327),
            .I(N__22082));
    ClkMux I__5287 (
            .O(N__22326),
            .I(N__22082));
    ClkMux I__5286 (
            .O(N__22325),
            .I(N__22082));
    ClkMux I__5285 (
            .O(N__22324),
            .I(N__22082));
    ClkMux I__5284 (
            .O(N__22323),
            .I(N__22082));
    ClkMux I__5283 (
            .O(N__22322),
            .I(N__22082));
    ClkMux I__5282 (
            .O(N__22321),
            .I(N__22082));
    ClkMux I__5281 (
            .O(N__22320),
            .I(N__22082));
    ClkMux I__5280 (
            .O(N__22319),
            .I(N__22082));
    ClkMux I__5279 (
            .O(N__22318),
            .I(N__22082));
    ClkMux I__5278 (
            .O(N__22317),
            .I(N__22082));
    ClkMux I__5277 (
            .O(N__22316),
            .I(N__22082));
    ClkMux I__5276 (
            .O(N__22315),
            .I(N__22082));
    ClkMux I__5275 (
            .O(N__22314),
            .I(N__22082));
    ClkMux I__5274 (
            .O(N__22313),
            .I(N__22082));
    ClkMux I__5273 (
            .O(N__22312),
            .I(N__22082));
    ClkMux I__5272 (
            .O(N__22311),
            .I(N__22082));
    ClkMux I__5271 (
            .O(N__22310),
            .I(N__22082));
    ClkMux I__5270 (
            .O(N__22309),
            .I(N__22082));
    ClkMux I__5269 (
            .O(N__22308),
            .I(N__22082));
    ClkMux I__5268 (
            .O(N__22307),
            .I(N__22082));
    ClkMux I__5267 (
            .O(N__22306),
            .I(N__22082));
    ClkMux I__5266 (
            .O(N__22305),
            .I(N__22082));
    ClkMux I__5265 (
            .O(N__22304),
            .I(N__22082));
    ClkMux I__5264 (
            .O(N__22303),
            .I(N__22082));
    ClkMux I__5263 (
            .O(N__22302),
            .I(N__22082));
    ClkMux I__5262 (
            .O(N__22301),
            .I(N__22082));
    ClkMux I__5261 (
            .O(N__22300),
            .I(N__22082));
    ClkMux I__5260 (
            .O(N__22299),
            .I(N__22082));
    ClkMux I__5259 (
            .O(N__22298),
            .I(N__22082));
    ClkMux I__5258 (
            .O(N__22297),
            .I(N__22082));
    ClkMux I__5257 (
            .O(N__22296),
            .I(N__22082));
    ClkMux I__5256 (
            .O(N__22295),
            .I(N__22082));
    ClkMux I__5255 (
            .O(N__22294),
            .I(N__22082));
    ClkMux I__5254 (
            .O(N__22293),
            .I(N__22082));
    ClkMux I__5253 (
            .O(N__22292),
            .I(N__22082));
    ClkMux I__5252 (
            .O(N__22291),
            .I(N__22082));
    ClkMux I__5251 (
            .O(N__22290),
            .I(N__22082));
    ClkMux I__5250 (
            .O(N__22289),
            .I(N__22082));
    ClkMux I__5249 (
            .O(N__22288),
            .I(N__22082));
    ClkMux I__5248 (
            .O(N__22287),
            .I(N__22082));
    ClkMux I__5247 (
            .O(N__22286),
            .I(N__22082));
    ClkMux I__5246 (
            .O(N__22285),
            .I(N__22082));
    ClkMux I__5245 (
            .O(N__22284),
            .I(N__22082));
    ClkMux I__5244 (
            .O(N__22283),
            .I(N__22082));
    ClkMux I__5243 (
            .O(N__22282),
            .I(N__22082));
    ClkMux I__5242 (
            .O(N__22281),
            .I(N__22082));
    ClkMux I__5241 (
            .O(N__22280),
            .I(N__22082));
    ClkMux I__5240 (
            .O(N__22279),
            .I(N__22082));
    ClkMux I__5239 (
            .O(N__22278),
            .I(N__22082));
    ClkMux I__5238 (
            .O(N__22277),
            .I(N__22082));
    ClkMux I__5237 (
            .O(N__22276),
            .I(N__22082));
    ClkMux I__5236 (
            .O(N__22275),
            .I(N__22082));
    ClkMux I__5235 (
            .O(N__22274),
            .I(N__22082));
    ClkMux I__5234 (
            .O(N__22273),
            .I(N__22082));
    ClkMux I__5233 (
            .O(N__22272),
            .I(N__22082));
    ClkMux I__5232 (
            .O(N__22271),
            .I(N__22082));
    ClkMux I__5231 (
            .O(N__22270),
            .I(N__22082));
    ClkMux I__5230 (
            .O(N__22269),
            .I(N__22082));
    GlobalMux I__5229 (
            .O(N__22082),
            .I(N__22079));
    gio2CtrlBuf I__5228 (
            .O(N__22079),
            .I(clk_g));
    CEMux I__5227 (
            .O(N__22076),
            .I(N__22046));
    CEMux I__5226 (
            .O(N__22075),
            .I(N__22046));
    CEMux I__5225 (
            .O(N__22074),
            .I(N__22046));
    CEMux I__5224 (
            .O(N__22073),
            .I(N__22046));
    CEMux I__5223 (
            .O(N__22072),
            .I(N__22046));
    CEMux I__5222 (
            .O(N__22071),
            .I(N__22046));
    CEMux I__5221 (
            .O(N__22070),
            .I(N__22046));
    CEMux I__5220 (
            .O(N__22069),
            .I(N__22046));
    CEMux I__5219 (
            .O(N__22068),
            .I(N__22046));
    CEMux I__5218 (
            .O(N__22067),
            .I(N__22046));
    GlobalMux I__5217 (
            .O(N__22046),
            .I(N__22043));
    gio2CtrlBuf I__5216 (
            .O(N__22043),
            .I(\buart.Z_rx.sample_g ));
    InMux I__5215 (
            .O(N__22040),
            .I(N__22031));
    InMux I__5214 (
            .O(N__22039),
            .I(N__22028));
    InMux I__5213 (
            .O(N__22038),
            .I(N__22025));
    InMux I__5212 (
            .O(N__22037),
            .I(N__22022));
    InMux I__5211 (
            .O(N__22036),
            .I(N__22019));
    SRMux I__5210 (
            .O(N__22035),
            .I(N__22014));
    InMux I__5209 (
            .O(N__22034),
            .I(N__22014));
    LocalMux I__5208 (
            .O(N__22031),
            .I(N__21966));
    LocalMux I__5207 (
            .O(N__22028),
            .I(N__21963));
    LocalMux I__5206 (
            .O(N__22025),
            .I(N__21960));
    LocalMux I__5205 (
            .O(N__22022),
            .I(N__21957));
    LocalMux I__5204 (
            .O(N__22019),
            .I(N__21954));
    LocalMux I__5203 (
            .O(N__22014),
            .I(N__21935));
    SRMux I__5202 (
            .O(N__22013),
            .I(N__21800));
    SRMux I__5201 (
            .O(N__22012),
            .I(N__21800));
    SRMux I__5200 (
            .O(N__22011),
            .I(N__21800));
    SRMux I__5199 (
            .O(N__22010),
            .I(N__21800));
    SRMux I__5198 (
            .O(N__22009),
            .I(N__21800));
    SRMux I__5197 (
            .O(N__22008),
            .I(N__21800));
    SRMux I__5196 (
            .O(N__22007),
            .I(N__21800));
    SRMux I__5195 (
            .O(N__22006),
            .I(N__21800));
    SRMux I__5194 (
            .O(N__22005),
            .I(N__21800));
    SRMux I__5193 (
            .O(N__22004),
            .I(N__21800));
    SRMux I__5192 (
            .O(N__22003),
            .I(N__21800));
    SRMux I__5191 (
            .O(N__22002),
            .I(N__21800));
    SRMux I__5190 (
            .O(N__22001),
            .I(N__21800));
    SRMux I__5189 (
            .O(N__22000),
            .I(N__21800));
    SRMux I__5188 (
            .O(N__21999),
            .I(N__21800));
    SRMux I__5187 (
            .O(N__21998),
            .I(N__21800));
    SRMux I__5186 (
            .O(N__21997),
            .I(N__21800));
    SRMux I__5185 (
            .O(N__21996),
            .I(N__21800));
    SRMux I__5184 (
            .O(N__21995),
            .I(N__21800));
    SRMux I__5183 (
            .O(N__21994),
            .I(N__21800));
    SRMux I__5182 (
            .O(N__21993),
            .I(N__21800));
    SRMux I__5181 (
            .O(N__21992),
            .I(N__21800));
    SRMux I__5180 (
            .O(N__21991),
            .I(N__21800));
    SRMux I__5179 (
            .O(N__21990),
            .I(N__21800));
    SRMux I__5178 (
            .O(N__21989),
            .I(N__21800));
    SRMux I__5177 (
            .O(N__21988),
            .I(N__21800));
    SRMux I__5176 (
            .O(N__21987),
            .I(N__21800));
    SRMux I__5175 (
            .O(N__21986),
            .I(N__21800));
    SRMux I__5174 (
            .O(N__21985),
            .I(N__21800));
    SRMux I__5173 (
            .O(N__21984),
            .I(N__21800));
    SRMux I__5172 (
            .O(N__21983),
            .I(N__21800));
    SRMux I__5171 (
            .O(N__21982),
            .I(N__21800));
    SRMux I__5170 (
            .O(N__21981),
            .I(N__21800));
    SRMux I__5169 (
            .O(N__21980),
            .I(N__21800));
    SRMux I__5168 (
            .O(N__21979),
            .I(N__21800));
    SRMux I__5167 (
            .O(N__21978),
            .I(N__21800));
    SRMux I__5166 (
            .O(N__21977),
            .I(N__21800));
    SRMux I__5165 (
            .O(N__21976),
            .I(N__21800));
    SRMux I__5164 (
            .O(N__21975),
            .I(N__21800));
    SRMux I__5163 (
            .O(N__21974),
            .I(N__21800));
    SRMux I__5162 (
            .O(N__21973),
            .I(N__21800));
    SRMux I__5161 (
            .O(N__21972),
            .I(N__21800));
    SRMux I__5160 (
            .O(N__21971),
            .I(N__21800));
    SRMux I__5159 (
            .O(N__21970),
            .I(N__21800));
    SRMux I__5158 (
            .O(N__21969),
            .I(N__21800));
    Glb2LocalMux I__5157 (
            .O(N__21966),
            .I(N__21800));
    Glb2LocalMux I__5156 (
            .O(N__21963),
            .I(N__21800));
    Glb2LocalMux I__5155 (
            .O(N__21960),
            .I(N__21800));
    Glb2LocalMux I__5154 (
            .O(N__21957),
            .I(N__21800));
    Glb2LocalMux I__5153 (
            .O(N__21954),
            .I(N__21800));
    SRMux I__5152 (
            .O(N__21953),
            .I(N__21800));
    SRMux I__5151 (
            .O(N__21952),
            .I(N__21800));
    SRMux I__5150 (
            .O(N__21951),
            .I(N__21800));
    SRMux I__5149 (
            .O(N__21950),
            .I(N__21800));
    SRMux I__5148 (
            .O(N__21949),
            .I(N__21800));
    SRMux I__5147 (
            .O(N__21948),
            .I(N__21800));
    SRMux I__5146 (
            .O(N__21947),
            .I(N__21800));
    SRMux I__5145 (
            .O(N__21946),
            .I(N__21800));
    SRMux I__5144 (
            .O(N__21945),
            .I(N__21800));
    SRMux I__5143 (
            .O(N__21944),
            .I(N__21800));
    SRMux I__5142 (
            .O(N__21943),
            .I(N__21800));
    SRMux I__5141 (
            .O(N__21942),
            .I(N__21800));
    SRMux I__5140 (
            .O(N__21941),
            .I(N__21800));
    SRMux I__5139 (
            .O(N__21940),
            .I(N__21800));
    SRMux I__5138 (
            .O(N__21939),
            .I(N__21800));
    SRMux I__5137 (
            .O(N__21938),
            .I(N__21800));
    Glb2LocalMux I__5136 (
            .O(N__21935),
            .I(N__21800));
    GlobalMux I__5135 (
            .O(N__21800),
            .I(N__21797));
    gio2CtrlBuf I__5134 (
            .O(N__21797),
            .I(rst_g));
    CascadeMux I__5133 (
            .O(N__21794),
            .I(N__21787));
    InMux I__5132 (
            .O(N__21793),
            .I(N__21781));
    CascadeMux I__5131 (
            .O(N__21792),
            .I(N__21778));
    CascadeMux I__5130 (
            .O(N__21791),
            .I(N__21769));
    CascadeMux I__5129 (
            .O(N__21790),
            .I(N__21765));
    InMux I__5128 (
            .O(N__21787),
            .I(N__21754));
    InMux I__5127 (
            .O(N__21786),
            .I(N__21754));
    InMux I__5126 (
            .O(N__21785),
            .I(N__21754));
    InMux I__5125 (
            .O(N__21784),
            .I(N__21754));
    LocalMux I__5124 (
            .O(N__21781),
            .I(N__21749));
    InMux I__5123 (
            .O(N__21778),
            .I(N__21746));
    InMux I__5122 (
            .O(N__21777),
            .I(N__21741));
    InMux I__5121 (
            .O(N__21776),
            .I(N__21741));
    InMux I__5120 (
            .O(N__21775),
            .I(N__21729));
    InMux I__5119 (
            .O(N__21774),
            .I(N__21729));
    InMux I__5118 (
            .O(N__21773),
            .I(N__21729));
    InMux I__5117 (
            .O(N__21772),
            .I(N__21729));
    InMux I__5116 (
            .O(N__21769),
            .I(N__21722));
    InMux I__5115 (
            .O(N__21768),
            .I(N__21722));
    InMux I__5114 (
            .O(N__21765),
            .I(N__21722));
    InMux I__5113 (
            .O(N__21764),
            .I(N__21719));
    CascadeMux I__5112 (
            .O(N__21763),
            .I(N__21714));
    LocalMux I__5111 (
            .O(N__21754),
            .I(N__21708));
    InMux I__5110 (
            .O(N__21753),
            .I(N__21705));
    CascadeMux I__5109 (
            .O(N__21752),
            .I(N__21702));
    Span4Mux_v I__5108 (
            .O(N__21749),
            .I(N__21699));
    LocalMux I__5107 (
            .O(N__21746),
            .I(N__21694));
    LocalMux I__5106 (
            .O(N__21741),
            .I(N__21694));
    InMux I__5105 (
            .O(N__21740),
            .I(N__21686));
    InMux I__5104 (
            .O(N__21739),
            .I(N__21686));
    InMux I__5103 (
            .O(N__21738),
            .I(N__21686));
    LocalMux I__5102 (
            .O(N__21729),
            .I(N__21679));
    LocalMux I__5101 (
            .O(N__21722),
            .I(N__21679));
    LocalMux I__5100 (
            .O(N__21719),
            .I(N__21679));
    InMux I__5099 (
            .O(N__21718),
            .I(N__21674));
    InMux I__5098 (
            .O(N__21717),
            .I(N__21674));
    InMux I__5097 (
            .O(N__21714),
            .I(N__21665));
    InMux I__5096 (
            .O(N__21713),
            .I(N__21665));
    InMux I__5095 (
            .O(N__21712),
            .I(N__21665));
    InMux I__5094 (
            .O(N__21711),
            .I(N__21665));
    Span4Mux_h I__5093 (
            .O(N__21708),
            .I(N__21662));
    LocalMux I__5092 (
            .O(N__21705),
            .I(N__21659));
    InMux I__5091 (
            .O(N__21702),
            .I(N__21656));
    Span4Mux_s3_h I__5090 (
            .O(N__21699),
            .I(N__21651));
    Span4Mux_v I__5089 (
            .O(N__21694),
            .I(N__21651));
    InMux I__5088 (
            .O(N__21693),
            .I(N__21648));
    LocalMux I__5087 (
            .O(N__21686),
            .I(N__21645));
    Span4Mux_v I__5086 (
            .O(N__21679),
            .I(N__21642));
    LocalMux I__5085 (
            .O(N__21674),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__5084 (
            .O(N__21665),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5083 (
            .O(N__21662),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5082 (
            .O(N__21659),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__5081 (
            .O(N__21656),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5080 (
            .O(N__21651),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__5079 (
            .O(N__21648),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5078 (
            .O(N__21645),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5077 (
            .O(N__21642),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    CascadeMux I__5076 (
            .O(N__21623),
            .I(\Lab_UT.dictrl.N_21_cascade_ ));
    InMux I__5075 (
            .O(N__21620),
            .I(N__21614));
    InMux I__5074 (
            .O(N__21619),
            .I(N__21614));
    LocalMux I__5073 (
            .O(N__21614),
            .I(N__21611));
    Span4Mux_h I__5072 (
            .O(N__21611),
            .I(N__21608));
    Odrv4 I__5071 (
            .O(N__21608),
            .I(\Lab_UT.dictrl.next_state_latmux_0_1 ));
    InMux I__5070 (
            .O(N__21605),
            .I(N__21598));
    InMux I__5069 (
            .O(N__21604),
            .I(N__21591));
    InMux I__5068 (
            .O(N__21603),
            .I(N__21591));
    InMux I__5067 (
            .O(N__21602),
            .I(N__21591));
    InMux I__5066 (
            .O(N__21601),
            .I(N__21588));
    LocalMux I__5065 (
            .O(N__21598),
            .I(N__21583));
    LocalMux I__5064 (
            .O(N__21591),
            .I(N__21583));
    LocalMux I__5063 (
            .O(N__21588),
            .I(N__21580));
    Span4Mux_v I__5062 (
            .O(N__21583),
            .I(N__21577));
    Odrv4 I__5061 (
            .O(N__21580),
            .I(\Lab_UT.dictrl.next_state18 ));
    Odrv4 I__5060 (
            .O(N__21577),
            .I(\Lab_UT.dictrl.next_state18 ));
    InMux I__5059 (
            .O(N__21572),
            .I(N__21565));
    CascadeMux I__5058 (
            .O(N__21571),
            .I(N__21561));
    InMux I__5057 (
            .O(N__21570),
            .I(N__21556));
    InMux I__5056 (
            .O(N__21569),
            .I(N__21556));
    InMux I__5055 (
            .O(N__21568),
            .I(N__21551));
    LocalMux I__5054 (
            .O(N__21565),
            .I(N__21548));
    InMux I__5053 (
            .O(N__21564),
            .I(N__21545));
    InMux I__5052 (
            .O(N__21561),
            .I(N__21542));
    LocalMux I__5051 (
            .O(N__21556),
            .I(N__21539));
    InMux I__5050 (
            .O(N__21555),
            .I(N__21536));
    CascadeMux I__5049 (
            .O(N__21554),
            .I(N__21531));
    LocalMux I__5048 (
            .O(N__21551),
            .I(N__21527));
    Span4Mux_h I__5047 (
            .O(N__21548),
            .I(N__21524));
    LocalMux I__5046 (
            .O(N__21545),
            .I(N__21519));
    LocalMux I__5045 (
            .O(N__21542),
            .I(N__21519));
    Span4Mux_h I__5044 (
            .O(N__21539),
            .I(N__21516));
    LocalMux I__5043 (
            .O(N__21536),
            .I(N__21513));
    InMux I__5042 (
            .O(N__21535),
            .I(N__21508));
    InMux I__5041 (
            .O(N__21534),
            .I(N__21508));
    InMux I__5040 (
            .O(N__21531),
            .I(N__21503));
    InMux I__5039 (
            .O(N__21530),
            .I(N__21503));
    Span4Mux_s2_h I__5038 (
            .O(N__21527),
            .I(N__21500));
    Odrv4 I__5037 (
            .O(N__21524),
            .I(bu_rx_data_1_rep2));
    Odrv12 I__5036 (
            .O(N__21519),
            .I(bu_rx_data_1_rep2));
    Odrv4 I__5035 (
            .O(N__21516),
            .I(bu_rx_data_1_rep2));
    Odrv4 I__5034 (
            .O(N__21513),
            .I(bu_rx_data_1_rep2));
    LocalMux I__5033 (
            .O(N__21508),
            .I(bu_rx_data_1_rep2));
    LocalMux I__5032 (
            .O(N__21503),
            .I(bu_rx_data_1_rep2));
    Odrv4 I__5031 (
            .O(N__21500),
            .I(bu_rx_data_1_rep2));
    CascadeMux I__5030 (
            .O(N__21485),
            .I(N__21482));
    InMux I__5029 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__5028 (
            .O(N__21479),
            .I(N__21476));
    Span4Mux_h I__5027 (
            .O(N__21476),
            .I(N__21473));
    Odrv4 I__5026 (
            .O(N__21473),
            .I(\Lab_UT.dictrl.g1_5_0 ));
    InMux I__5025 (
            .O(N__21470),
            .I(N__21456));
    InMux I__5024 (
            .O(N__21469),
            .I(N__21456));
    InMux I__5023 (
            .O(N__21468),
            .I(N__21456));
    InMux I__5022 (
            .O(N__21467),
            .I(N__21456));
    CascadeMux I__5021 (
            .O(N__21466),
            .I(N__21449));
    InMux I__5020 (
            .O(N__21465),
            .I(N__21443));
    LocalMux I__5019 (
            .O(N__21456),
            .I(N__21440));
    InMux I__5018 (
            .O(N__21455),
            .I(N__21435));
    InMux I__5017 (
            .O(N__21454),
            .I(N__21435));
    InMux I__5016 (
            .O(N__21453),
            .I(N__21424));
    InMux I__5015 (
            .O(N__21452),
            .I(N__21420));
    InMux I__5014 (
            .O(N__21449),
            .I(N__21411));
    InMux I__5013 (
            .O(N__21448),
            .I(N__21411));
    InMux I__5012 (
            .O(N__21447),
            .I(N__21411));
    InMux I__5011 (
            .O(N__21446),
            .I(N__21411));
    LocalMux I__5010 (
            .O(N__21443),
            .I(N__21406));
    Span4Mux_v I__5009 (
            .O(N__21440),
            .I(N__21406));
    LocalMux I__5008 (
            .O(N__21435),
            .I(N__21403));
    InMux I__5007 (
            .O(N__21434),
            .I(N__21400));
    CascadeMux I__5006 (
            .O(N__21433),
            .I(N__21397));
    InMux I__5005 (
            .O(N__21432),
            .I(N__21392));
    InMux I__5004 (
            .O(N__21431),
            .I(N__21392));
    InMux I__5003 (
            .O(N__21430),
            .I(N__21387));
    InMux I__5002 (
            .O(N__21429),
            .I(N__21387));
    InMux I__5001 (
            .O(N__21428),
            .I(N__21384));
    InMux I__5000 (
            .O(N__21427),
            .I(N__21381));
    LocalMux I__4999 (
            .O(N__21424),
            .I(N__21378));
    CascadeMux I__4998 (
            .O(N__21423),
            .I(N__21370));
    LocalMux I__4997 (
            .O(N__21420),
            .I(N__21366));
    LocalMux I__4996 (
            .O(N__21411),
            .I(N__21356));
    Span4Mux_h I__4995 (
            .O(N__21406),
            .I(N__21356));
    Span4Mux_v I__4994 (
            .O(N__21403),
            .I(N__21356));
    LocalMux I__4993 (
            .O(N__21400),
            .I(N__21353));
    InMux I__4992 (
            .O(N__21397),
            .I(N__21350));
    LocalMux I__4991 (
            .O(N__21392),
            .I(N__21347));
    LocalMux I__4990 (
            .O(N__21387),
            .I(N__21340));
    LocalMux I__4989 (
            .O(N__21384),
            .I(N__21340));
    LocalMux I__4988 (
            .O(N__21381),
            .I(N__21340));
    Span4Mux_h I__4987 (
            .O(N__21378),
            .I(N__21337));
    InMux I__4986 (
            .O(N__21377),
            .I(N__21334));
    InMux I__4985 (
            .O(N__21376),
            .I(N__21323));
    InMux I__4984 (
            .O(N__21375),
            .I(N__21323));
    InMux I__4983 (
            .O(N__21374),
            .I(N__21323));
    InMux I__4982 (
            .O(N__21373),
            .I(N__21323));
    InMux I__4981 (
            .O(N__21370),
            .I(N__21323));
    InMux I__4980 (
            .O(N__21369),
            .I(N__21320));
    Span4Mux_h I__4979 (
            .O(N__21366),
            .I(N__21317));
    InMux I__4978 (
            .O(N__21365),
            .I(N__21310));
    InMux I__4977 (
            .O(N__21364),
            .I(N__21310));
    InMux I__4976 (
            .O(N__21363),
            .I(N__21310));
    Sp12to4 I__4975 (
            .O(N__21356),
            .I(N__21307));
    Span4Mux_s3_h I__4974 (
            .O(N__21353),
            .I(N__21296));
    LocalMux I__4973 (
            .O(N__21350),
            .I(N__21296));
    Span4Mux_h I__4972 (
            .O(N__21347),
            .I(N__21296));
    Span4Mux_h I__4971 (
            .O(N__21340),
            .I(N__21296));
    Span4Mux_h I__4970 (
            .O(N__21337),
            .I(N__21296));
    LocalMux I__4969 (
            .O(N__21334),
            .I(\Lab_UT.state_1 ));
    LocalMux I__4968 (
            .O(N__21323),
            .I(\Lab_UT.state_1 ));
    LocalMux I__4967 (
            .O(N__21320),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__4966 (
            .O(N__21317),
            .I(\Lab_UT.state_1 ));
    LocalMux I__4965 (
            .O(N__21310),
            .I(\Lab_UT.state_1 ));
    Odrv12 I__4964 (
            .O(N__21307),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__4963 (
            .O(N__21296),
            .I(\Lab_UT.state_1 ));
    InMux I__4962 (
            .O(N__21281),
            .I(N__21277));
    InMux I__4961 (
            .O(N__21280),
            .I(N__21274));
    LocalMux I__4960 (
            .O(N__21277),
            .I(\Lab_UT.dictrl.N_23 ));
    LocalMux I__4959 (
            .O(N__21274),
            .I(\Lab_UT.dictrl.N_23 ));
    InMux I__4958 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__4957 (
            .O(N__21266),
            .I(N__21263));
    Span4Mux_h I__4956 (
            .O(N__21263),
            .I(N__21260));
    Odrv4 I__4955 (
            .O(N__21260),
            .I(\Lab_UT.dictrl.N_30 ));
    CascadeMux I__4954 (
            .O(N__21257),
            .I(\Lab_UT.dictrl.next_state5_3_cascade_ ));
    InMux I__4953 (
            .O(N__21254),
            .I(N__21251));
    LocalMux I__4952 (
            .O(N__21251),
            .I(N__21248));
    Span4Mux_s2_h I__4951 (
            .O(N__21248),
            .I(N__21244));
    InMux I__4950 (
            .O(N__21247),
            .I(N__21241));
    Odrv4 I__4949 (
            .O(N__21244),
            .I(\Lab_UT.dictrl.next_state32Z0Z_1 ));
    LocalMux I__4948 (
            .O(N__21241),
            .I(\Lab_UT.dictrl.next_state32Z0Z_1 ));
    CascadeMux I__4947 (
            .O(N__21236),
            .I(N__21232));
    CascadeMux I__4946 (
            .O(N__21235),
            .I(N__21229));
    InMux I__4945 (
            .O(N__21232),
            .I(N__21224));
    InMux I__4944 (
            .O(N__21229),
            .I(N__21224));
    LocalMux I__4943 (
            .O(N__21224),
            .I(N__21221));
    Span4Mux_h I__4942 (
            .O(N__21221),
            .I(N__21218));
    Sp12to4 I__4941 (
            .O(N__21218),
            .I(N__21215));
    Odrv12 I__4940 (
            .O(N__21215),
            .I(\Lab_UT.dictrl.N_18 ));
    InMux I__4939 (
            .O(N__21212),
            .I(N__21203));
    InMux I__4938 (
            .O(N__21211),
            .I(N__21203));
    InMux I__4937 (
            .O(N__21210),
            .I(N__21199));
    InMux I__4936 (
            .O(N__21209),
            .I(N__21195));
    InMux I__4935 (
            .O(N__21208),
            .I(N__21192));
    LocalMux I__4934 (
            .O(N__21203),
            .I(N__21189));
    InMux I__4933 (
            .O(N__21202),
            .I(N__21186));
    LocalMux I__4932 (
            .O(N__21199),
            .I(N__21183));
    CascadeMux I__4931 (
            .O(N__21198),
            .I(N__21179));
    LocalMux I__4930 (
            .O(N__21195),
            .I(N__21174));
    LocalMux I__4929 (
            .O(N__21192),
            .I(N__21174));
    Span4Mux_v I__4928 (
            .O(N__21189),
            .I(N__21169));
    LocalMux I__4927 (
            .O(N__21186),
            .I(N__21169));
    Span4Mux_h I__4926 (
            .O(N__21183),
            .I(N__21166));
    InMux I__4925 (
            .O(N__21182),
            .I(N__21163));
    InMux I__4924 (
            .O(N__21179),
            .I(N__21160));
    Span4Mux_v I__4923 (
            .O(N__21174),
            .I(N__21157));
    Span4Mux_h I__4922 (
            .O(N__21169),
            .I(N__21154));
    Sp12to4 I__4921 (
            .O(N__21166),
            .I(N__21147));
    LocalMux I__4920 (
            .O(N__21163),
            .I(N__21147));
    LocalMux I__4919 (
            .O(N__21160),
            .I(N__21147));
    Odrv4 I__4918 (
            .O(N__21157),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    Odrv4 I__4917 (
            .O(N__21154),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    Odrv12 I__4916 (
            .O(N__21147),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    InMux I__4915 (
            .O(N__21140),
            .I(N__21137));
    LocalMux I__4914 (
            .O(N__21137),
            .I(\Lab_UT.dictrl.m17_1 ));
    InMux I__4913 (
            .O(N__21134),
            .I(N__21118));
    InMux I__4912 (
            .O(N__21133),
            .I(N__21118));
    CascadeMux I__4911 (
            .O(N__21132),
            .I(N__21115));
    InMux I__4910 (
            .O(N__21131),
            .I(N__21105));
    InMux I__4909 (
            .O(N__21130),
            .I(N__21100));
    InMux I__4908 (
            .O(N__21129),
            .I(N__21100));
    InMux I__4907 (
            .O(N__21128),
            .I(N__21095));
    InMux I__4906 (
            .O(N__21127),
            .I(N__21095));
    InMux I__4905 (
            .O(N__21126),
            .I(N__21092));
    InMux I__4904 (
            .O(N__21125),
            .I(N__21087));
    InMux I__4903 (
            .O(N__21124),
            .I(N__21087));
    InMux I__4902 (
            .O(N__21123),
            .I(N__21084));
    LocalMux I__4901 (
            .O(N__21118),
            .I(N__21081));
    InMux I__4900 (
            .O(N__21115),
            .I(N__21074));
    InMux I__4899 (
            .O(N__21114),
            .I(N__21074));
    InMux I__4898 (
            .O(N__21113),
            .I(N__21074));
    InMux I__4897 (
            .O(N__21112),
            .I(N__21068));
    InMux I__4896 (
            .O(N__21111),
            .I(N__21056));
    InMux I__4895 (
            .O(N__21110),
            .I(N__21051));
    InMux I__4894 (
            .O(N__21109),
            .I(N__21051));
    InMux I__4893 (
            .O(N__21108),
            .I(N__21048));
    LocalMux I__4892 (
            .O(N__21105),
            .I(N__21043));
    LocalMux I__4891 (
            .O(N__21100),
            .I(N__21043));
    LocalMux I__4890 (
            .O(N__21095),
            .I(N__21036));
    LocalMux I__4889 (
            .O(N__21092),
            .I(N__21036));
    LocalMux I__4888 (
            .O(N__21087),
            .I(N__21036));
    LocalMux I__4887 (
            .O(N__21084),
            .I(N__21033));
    Span4Mux_v I__4886 (
            .O(N__21081),
            .I(N__21028));
    LocalMux I__4885 (
            .O(N__21074),
            .I(N__21028));
    InMux I__4884 (
            .O(N__21073),
            .I(N__21023));
    InMux I__4883 (
            .O(N__21072),
            .I(N__21023));
    InMux I__4882 (
            .O(N__21071),
            .I(N__21020));
    LocalMux I__4881 (
            .O(N__21068),
            .I(N__21017));
    InMux I__4880 (
            .O(N__21067),
            .I(N__21010));
    InMux I__4879 (
            .O(N__21066),
            .I(N__21010));
    InMux I__4878 (
            .O(N__21065),
            .I(N__21010));
    InMux I__4877 (
            .O(N__21064),
            .I(N__21007));
    InMux I__4876 (
            .O(N__21063),
            .I(N__21002));
    InMux I__4875 (
            .O(N__21062),
            .I(N__21002));
    InMux I__4874 (
            .O(N__21061),
            .I(N__20995));
    InMux I__4873 (
            .O(N__21060),
            .I(N__20995));
    InMux I__4872 (
            .O(N__21059),
            .I(N__20995));
    LocalMux I__4871 (
            .O(N__21056),
            .I(N__20988));
    LocalMux I__4870 (
            .O(N__21051),
            .I(N__20988));
    LocalMux I__4869 (
            .O(N__21048),
            .I(N__20988));
    Span4Mux_v I__4868 (
            .O(N__21043),
            .I(N__20983));
    Span4Mux_v I__4867 (
            .O(N__21036),
            .I(N__20983));
    Span4Mux_v I__4866 (
            .O(N__21033),
            .I(N__20980));
    Span4Mux_s3_h I__4865 (
            .O(N__21028),
            .I(N__20977));
    LocalMux I__4864 (
            .O(N__21023),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4863 (
            .O(N__21020),
            .I(\Lab_UT.state_0 ));
    Odrv12 I__4862 (
            .O(N__21017),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4861 (
            .O(N__21010),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4860 (
            .O(N__21007),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4859 (
            .O(N__21002),
            .I(\Lab_UT.state_0 ));
    LocalMux I__4858 (
            .O(N__20995),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__4857 (
            .O(N__20988),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__4856 (
            .O(N__20983),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__4855 (
            .O(N__20980),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__4854 (
            .O(N__20977),
            .I(\Lab_UT.state_0 ));
    InMux I__4853 (
            .O(N__20954),
            .I(N__20944));
    InMux I__4852 (
            .O(N__20953),
            .I(N__20944));
    InMux I__4851 (
            .O(N__20952),
            .I(N__20936));
    InMux I__4850 (
            .O(N__20951),
            .I(N__20936));
    InMux I__4849 (
            .O(N__20950),
            .I(N__20936));
    InMux I__4848 (
            .O(N__20949),
            .I(N__20933));
    LocalMux I__4847 (
            .O(N__20944),
            .I(N__20930));
    InMux I__4846 (
            .O(N__20943),
            .I(N__20927));
    LocalMux I__4845 (
            .O(N__20936),
            .I(N__20924));
    LocalMux I__4844 (
            .O(N__20933),
            .I(N__20921));
    Span4Mux_s2_h I__4843 (
            .O(N__20930),
            .I(N__20918));
    LocalMux I__4842 (
            .O(N__20927),
            .I(\Lab_UT.dictrl.next_stateZ0Z32 ));
    Odrv12 I__4841 (
            .O(N__20924),
            .I(\Lab_UT.dictrl.next_stateZ0Z32 ));
    Odrv4 I__4840 (
            .O(N__20921),
            .I(\Lab_UT.dictrl.next_stateZ0Z32 ));
    Odrv4 I__4839 (
            .O(N__20918),
            .I(\Lab_UT.dictrl.next_stateZ0Z32 ));
    InMux I__4838 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__4837 (
            .O(N__20906),
            .I(\Lab_UT.dictrl.N_29_0 ));
    CascadeMux I__4836 (
            .O(N__20903),
            .I(N__20900));
    InMux I__4835 (
            .O(N__20900),
            .I(N__20896));
    CascadeMux I__4834 (
            .O(N__20899),
            .I(N__20893));
    LocalMux I__4833 (
            .O(N__20896),
            .I(N__20890));
    InMux I__4832 (
            .O(N__20893),
            .I(N__20887));
    Span4Mux_h I__4831 (
            .O(N__20890),
            .I(N__20882));
    LocalMux I__4830 (
            .O(N__20887),
            .I(N__20882));
    Span4Mux_s2_h I__4829 (
            .O(N__20882),
            .I(N__20879));
    Odrv4 I__4828 (
            .O(N__20879),
            .I(bu_rx_data_fast_0));
    InMux I__4827 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__4826 (
            .O(N__20873),
            .I(N__20870));
    Odrv4 I__4825 (
            .O(N__20870),
            .I(\Lab_UT.dictrl.g0_0_0_a3_1 ));
    CascadeMux I__4824 (
            .O(N__20867),
            .I(N__20862));
    CascadeMux I__4823 (
            .O(N__20866),
            .I(N__20859));
    InMux I__4822 (
            .O(N__20865),
            .I(N__20833));
    InMux I__4821 (
            .O(N__20862),
            .I(N__20833));
    InMux I__4820 (
            .O(N__20859),
            .I(N__20833));
    InMux I__4819 (
            .O(N__20858),
            .I(N__20833));
    InMux I__4818 (
            .O(N__20857),
            .I(N__20833));
    InMux I__4817 (
            .O(N__20856),
            .I(N__20833));
    InMux I__4816 (
            .O(N__20855),
            .I(N__20833));
    CascadeMux I__4815 (
            .O(N__20854),
            .I(N__20830));
    InMux I__4814 (
            .O(N__20853),
            .I(N__20825));
    InMux I__4813 (
            .O(N__20852),
            .I(N__20818));
    InMux I__4812 (
            .O(N__20851),
            .I(N__20818));
    InMux I__4811 (
            .O(N__20850),
            .I(N__20818));
    InMux I__4810 (
            .O(N__20849),
            .I(N__20812));
    InMux I__4809 (
            .O(N__20848),
            .I(N__20812));
    LocalMux I__4808 (
            .O(N__20833),
            .I(N__20808));
    InMux I__4807 (
            .O(N__20830),
            .I(N__20801));
    InMux I__4806 (
            .O(N__20829),
            .I(N__20801));
    InMux I__4805 (
            .O(N__20828),
            .I(N__20801));
    LocalMux I__4804 (
            .O(N__20825),
            .I(N__20790));
    LocalMux I__4803 (
            .O(N__20818),
            .I(N__20790));
    InMux I__4802 (
            .O(N__20817),
            .I(N__20787));
    LocalMux I__4801 (
            .O(N__20812),
            .I(N__20784));
    InMux I__4800 (
            .O(N__20811),
            .I(N__20781));
    Span4Mux_v I__4799 (
            .O(N__20808),
            .I(N__20778));
    LocalMux I__4798 (
            .O(N__20801),
            .I(N__20775));
    InMux I__4797 (
            .O(N__20800),
            .I(N__20764));
    InMux I__4796 (
            .O(N__20799),
            .I(N__20764));
    InMux I__4795 (
            .O(N__20798),
            .I(N__20764));
    InMux I__4794 (
            .O(N__20797),
            .I(N__20764));
    InMux I__4793 (
            .O(N__20796),
            .I(N__20764));
    InMux I__4792 (
            .O(N__20795),
            .I(N__20761));
    Span4Mux_h I__4791 (
            .O(N__20790),
            .I(N__20756));
    LocalMux I__4790 (
            .O(N__20787),
            .I(N__20756));
    Odrv4 I__4789 (
            .O(N__20784),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__4788 (
            .O(N__20781),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__4787 (
            .O(N__20778),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__4786 (
            .O(N__20775),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__4785 (
            .O(N__20764),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__4784 (
            .O(N__20761),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__4783 (
            .O(N__20756),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    InMux I__4782 (
            .O(N__20741),
            .I(N__20738));
    LocalMux I__4781 (
            .O(N__20738),
            .I(N__20735));
    Odrv12 I__4780 (
            .O(N__20735),
            .I(\Lab_UT.dictrl.g0_0_i_a3_1 ));
    InMux I__4779 (
            .O(N__20732),
            .I(N__20729));
    LocalMux I__4778 (
            .O(N__20729),
            .I(N__20722));
    InMux I__4777 (
            .O(N__20728),
            .I(N__20719));
    InMux I__4776 (
            .O(N__20727),
            .I(N__20716));
    InMux I__4775 (
            .O(N__20726),
            .I(N__20711));
    InMux I__4774 (
            .O(N__20725),
            .I(N__20711));
    Span4Mux_v I__4773 (
            .O(N__20722),
            .I(N__20708));
    LocalMux I__4772 (
            .O(N__20719),
            .I(N__20705));
    LocalMux I__4771 (
            .O(N__20716),
            .I(N__20698));
    LocalMux I__4770 (
            .O(N__20711),
            .I(N__20698));
    Span4Mux_h I__4769 (
            .O(N__20708),
            .I(N__20698));
    Span12Mux_s8_v I__4768 (
            .O(N__20705),
            .I(N__20695));
    Odrv4 I__4767 (
            .O(N__20698),
            .I(\Lab_UT.dicLdAStens_0 ));
    Odrv12 I__4766 (
            .O(N__20695),
            .I(\Lab_UT.dicLdAStens_0 ));
    CascadeMux I__4765 (
            .O(N__20690),
            .I(N__20686));
    CascadeMux I__4764 (
            .O(N__20689),
            .I(N__20683));
    InMux I__4763 (
            .O(N__20686),
            .I(N__20672));
    InMux I__4762 (
            .O(N__20683),
            .I(N__20672));
    InMux I__4761 (
            .O(N__20682),
            .I(N__20672));
    InMux I__4760 (
            .O(N__20681),
            .I(N__20672));
    LocalMux I__4759 (
            .O(N__20672),
            .I(N__20669));
    Odrv4 I__4758 (
            .O(N__20669),
            .I(\Lab_UT.dictrl.N_40_mux ));
    CascadeMux I__4757 (
            .O(N__20666),
            .I(N__20659));
    CascadeMux I__4756 (
            .O(N__20665),
            .I(N__20651));
    CascadeMux I__4755 (
            .O(N__20664),
            .I(N__20646));
    InMux I__4754 (
            .O(N__20663),
            .I(N__20642));
    CascadeMux I__4753 (
            .O(N__20662),
            .I(N__20639));
    InMux I__4752 (
            .O(N__20659),
            .I(N__20628));
    InMux I__4751 (
            .O(N__20658),
            .I(N__20628));
    InMux I__4750 (
            .O(N__20657),
            .I(N__20628));
    InMux I__4749 (
            .O(N__20656),
            .I(N__20628));
    InMux I__4748 (
            .O(N__20655),
            .I(N__20628));
    InMux I__4747 (
            .O(N__20654),
            .I(N__20623));
    InMux I__4746 (
            .O(N__20651),
            .I(N__20623));
    InMux I__4745 (
            .O(N__20650),
            .I(N__20620));
    InMux I__4744 (
            .O(N__20649),
            .I(N__20615));
    InMux I__4743 (
            .O(N__20646),
            .I(N__20615));
    InMux I__4742 (
            .O(N__20645),
            .I(N__20612));
    LocalMux I__4741 (
            .O(N__20642),
            .I(N__20609));
    InMux I__4740 (
            .O(N__20639),
            .I(N__20598));
    LocalMux I__4739 (
            .O(N__20628),
            .I(N__20591));
    LocalMux I__4738 (
            .O(N__20623),
            .I(N__20591));
    LocalMux I__4737 (
            .O(N__20620),
            .I(N__20591));
    LocalMux I__4736 (
            .O(N__20615),
            .I(N__20586));
    LocalMux I__4735 (
            .O(N__20612),
            .I(N__20586));
    Span4Mux_h I__4734 (
            .O(N__20609),
            .I(N__20583));
    InMux I__4733 (
            .O(N__20608),
            .I(N__20578));
    InMux I__4732 (
            .O(N__20607),
            .I(N__20578));
    InMux I__4731 (
            .O(N__20606),
            .I(N__20573));
    InMux I__4730 (
            .O(N__20605),
            .I(N__20573));
    InMux I__4729 (
            .O(N__20604),
            .I(N__20570));
    InMux I__4728 (
            .O(N__20603),
            .I(N__20563));
    InMux I__4727 (
            .O(N__20602),
            .I(N__20563));
    InMux I__4726 (
            .O(N__20601),
            .I(N__20563));
    LocalMux I__4725 (
            .O(N__20598),
            .I(N__20560));
    Span12Mux_s10_h I__4724 (
            .O(N__20591),
            .I(N__20557));
    Span4Mux_v I__4723 (
            .O(N__20586),
            .I(N__20548));
    Span4Mux_v I__4722 (
            .O(N__20583),
            .I(N__20548));
    LocalMux I__4721 (
            .O(N__20578),
            .I(N__20548));
    LocalMux I__4720 (
            .O(N__20573),
            .I(N__20548));
    LocalMux I__4719 (
            .O(N__20570),
            .I(\Lab_UT.state_3 ));
    LocalMux I__4718 (
            .O(N__20563),
            .I(\Lab_UT.state_3 ));
    Odrv12 I__4717 (
            .O(N__20560),
            .I(\Lab_UT.state_3 ));
    Odrv12 I__4716 (
            .O(N__20557),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__4715 (
            .O(N__20548),
            .I(\Lab_UT.state_3 ));
    CascadeMux I__4714 (
            .O(N__20537),
            .I(\Lab_UT.dictrl.N_13_cascade_ ));
    CascadeMux I__4713 (
            .O(N__20534),
            .I(N__20531));
    InMux I__4712 (
            .O(N__20531),
            .I(N__20528));
    LocalMux I__4711 (
            .O(N__20528),
            .I(N__20525));
    Span4Mux_h I__4710 (
            .O(N__20525),
            .I(N__20522));
    Odrv4 I__4709 (
            .O(N__20522),
            .I(\Lab_UT.dictrl.N_16 ));
    InMux I__4708 (
            .O(N__20519),
            .I(N__20516));
    LocalMux I__4707 (
            .O(N__20516),
            .I(N__20513));
    Span4Mux_v I__4706 (
            .O(N__20513),
            .I(N__20509));
    InMux I__4705 (
            .O(N__20512),
            .I(N__20506));
    Span4Mux_h I__4704 (
            .O(N__20509),
            .I(N__20501));
    LocalMux I__4703 (
            .O(N__20506),
            .I(N__20501));
    Odrv4 I__4702 (
            .O(N__20501),
            .I(\Lab_UT.dictrl.state_fast_3 ));
    CascadeMux I__4701 (
            .O(N__20498),
            .I(N__20495));
    InMux I__4700 (
            .O(N__20495),
            .I(N__20486));
    InMux I__4699 (
            .O(N__20494),
            .I(N__20486));
    CascadeMux I__4698 (
            .O(N__20493),
            .I(N__20483));
    InMux I__4697 (
            .O(N__20492),
            .I(N__20478));
    InMux I__4696 (
            .O(N__20491),
            .I(N__20475));
    LocalMux I__4695 (
            .O(N__20486),
            .I(N__20472));
    InMux I__4694 (
            .O(N__20483),
            .I(N__20469));
    InMux I__4693 (
            .O(N__20482),
            .I(N__20464));
    InMux I__4692 (
            .O(N__20481),
            .I(N__20464));
    LocalMux I__4691 (
            .O(N__20478),
            .I(N__20457));
    LocalMux I__4690 (
            .O(N__20475),
            .I(N__20454));
    Span4Mux_h I__4689 (
            .O(N__20472),
            .I(N__20451));
    LocalMux I__4688 (
            .O(N__20469),
            .I(N__20446));
    LocalMux I__4687 (
            .O(N__20464),
            .I(N__20446));
    InMux I__4686 (
            .O(N__20463),
            .I(N__20441));
    InMux I__4685 (
            .O(N__20462),
            .I(N__20441));
    InMux I__4684 (
            .O(N__20461),
            .I(N__20436));
    InMux I__4683 (
            .O(N__20460),
            .I(N__20436));
    Span4Mux_s2_h I__4682 (
            .O(N__20457),
            .I(N__20433));
    Odrv4 I__4681 (
            .O(N__20454),
            .I(bu_rx_data_2_rep2));
    Odrv4 I__4680 (
            .O(N__20451),
            .I(bu_rx_data_2_rep2));
    Odrv4 I__4679 (
            .O(N__20446),
            .I(bu_rx_data_2_rep2));
    LocalMux I__4678 (
            .O(N__20441),
            .I(bu_rx_data_2_rep2));
    LocalMux I__4677 (
            .O(N__20436),
            .I(bu_rx_data_2_rep2));
    Odrv4 I__4676 (
            .O(N__20433),
            .I(bu_rx_data_2_rep2));
    InMux I__4675 (
            .O(N__20420),
            .I(N__20417));
    LocalMux I__4674 (
            .O(N__20417),
            .I(\Lab_UT.dictrl.N_15 ));
    InMux I__4673 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__4672 (
            .O(N__20411),
            .I(N__20405));
    InMux I__4671 (
            .O(N__20410),
            .I(N__20402));
    InMux I__4670 (
            .O(N__20409),
            .I(N__20399));
    InMux I__4669 (
            .O(N__20408),
            .I(N__20396));
    Span4Mux_v I__4668 (
            .O(N__20405),
            .I(N__20391));
    LocalMux I__4667 (
            .O(N__20402),
            .I(N__20384));
    LocalMux I__4666 (
            .O(N__20399),
            .I(N__20384));
    LocalMux I__4665 (
            .O(N__20396),
            .I(N__20384));
    InMux I__4664 (
            .O(N__20395),
            .I(N__20381));
    InMux I__4663 (
            .O(N__20394),
            .I(N__20378));
    Span4Mux_h I__4662 (
            .O(N__20391),
            .I(N__20373));
    Span4Mux_s3_h I__4661 (
            .O(N__20384),
            .I(N__20373));
    LocalMux I__4660 (
            .O(N__20381),
            .I(N__20368));
    LocalMux I__4659 (
            .O(N__20378),
            .I(N__20368));
    Odrv4 I__4658 (
            .O(N__20373),
            .I(\Lab_UT.dictrl.next_state12 ));
    Odrv4 I__4657 (
            .O(N__20368),
            .I(\Lab_UT.dictrl.next_state12 ));
    InMux I__4656 (
            .O(N__20363),
            .I(N__20360));
    LocalMux I__4655 (
            .O(N__20360),
            .I(N__20357));
    Odrv4 I__4654 (
            .O(N__20357),
            .I(\Lab_UT.bcd2segment4.segment_0Z0Z_0 ));
    InMux I__4653 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__4652 (
            .O(N__20351),
            .I(N__20348));
    Odrv4 I__4651 (
            .O(N__20348),
            .I(\Lab_UT.bcd2segment4.segment_0Z0Z_1 ));
    CascadeMux I__4650 (
            .O(N__20345),
            .I(N__20335));
    InMux I__4649 (
            .O(N__20344),
            .I(N__20320));
    InMux I__4648 (
            .O(N__20343),
            .I(N__20320));
    InMux I__4647 (
            .O(N__20342),
            .I(N__20320));
    InMux I__4646 (
            .O(N__20341),
            .I(N__20320));
    InMux I__4645 (
            .O(N__20340),
            .I(N__20320));
    InMux I__4644 (
            .O(N__20339),
            .I(N__20320));
    InMux I__4643 (
            .O(N__20338),
            .I(N__20320));
    InMux I__4642 (
            .O(N__20335),
            .I(N__20317));
    LocalMux I__4641 (
            .O(N__20320),
            .I(N__20313));
    LocalMux I__4640 (
            .O(N__20317),
            .I(N__20307));
    InMux I__4639 (
            .O(N__20316),
            .I(N__20304));
    Span4Mux_s3_h I__4638 (
            .O(N__20313),
            .I(N__20301));
    InMux I__4637 (
            .O(N__20312),
            .I(N__20298));
    InMux I__4636 (
            .O(N__20311),
            .I(N__20293));
    InMux I__4635 (
            .O(N__20310),
            .I(N__20293));
    Span4Mux_h I__4634 (
            .O(N__20307),
            .I(N__20290));
    LocalMux I__4633 (
            .O(N__20304),
            .I(N__20285));
    Span4Mux_v I__4632 (
            .O(N__20301),
            .I(N__20285));
    LocalMux I__4631 (
            .O(N__20298),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__4630 (
            .O(N__20293),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__4629 (
            .O(N__20290),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__4628 (
            .O(N__20285),
            .I(\Lab_UT.di_Mtens_2 ));
    CascadeMux I__4627 (
            .O(N__20276),
            .I(N__20269));
    CascadeMux I__4626 (
            .O(N__20275),
            .I(N__20265));
    CascadeMux I__4625 (
            .O(N__20274),
            .I(N__20261));
    InMux I__4624 (
            .O(N__20273),
            .I(N__20246));
    InMux I__4623 (
            .O(N__20272),
            .I(N__20246));
    InMux I__4622 (
            .O(N__20269),
            .I(N__20246));
    InMux I__4621 (
            .O(N__20268),
            .I(N__20246));
    InMux I__4620 (
            .O(N__20265),
            .I(N__20246));
    InMux I__4619 (
            .O(N__20264),
            .I(N__20246));
    InMux I__4618 (
            .O(N__20261),
            .I(N__20246));
    LocalMux I__4617 (
            .O(N__20246),
            .I(N__20243));
    Span4Mux_s1_h I__4616 (
            .O(N__20243),
            .I(N__20237));
    InMux I__4615 (
            .O(N__20242),
            .I(N__20234));
    InMux I__4614 (
            .O(N__20241),
            .I(N__20229));
    InMux I__4613 (
            .O(N__20240),
            .I(N__20229));
    Span4Mux_h I__4612 (
            .O(N__20237),
            .I(N__20226));
    LocalMux I__4611 (
            .O(N__20234),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__4610 (
            .O(N__20229),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__4609 (
            .O(N__20226),
            .I(\Lab_UT.di_Mtens_3 ));
    CascadeMux I__4608 (
            .O(N__20219),
            .I(N__20210));
    CascadeMux I__4607 (
            .O(N__20218),
            .I(N__20207));
    CascadeMux I__4606 (
            .O(N__20217),
            .I(N__20204));
    CascadeMux I__4605 (
            .O(N__20216),
            .I(N__20201));
    InMux I__4604 (
            .O(N__20215),
            .I(N__20194));
    InMux I__4603 (
            .O(N__20214),
            .I(N__20194));
    InMux I__4602 (
            .O(N__20213),
            .I(N__20194));
    InMux I__4601 (
            .O(N__20210),
            .I(N__20185));
    InMux I__4600 (
            .O(N__20207),
            .I(N__20185));
    InMux I__4599 (
            .O(N__20204),
            .I(N__20185));
    InMux I__4598 (
            .O(N__20201),
            .I(N__20185));
    LocalMux I__4597 (
            .O(N__20194),
            .I(N__20179));
    LocalMux I__4596 (
            .O(N__20185),
            .I(N__20179));
    CascadeMux I__4595 (
            .O(N__20184),
            .I(N__20174));
    Span4Mux_s1_h I__4594 (
            .O(N__20179),
            .I(N__20169));
    InMux I__4593 (
            .O(N__20178),
            .I(N__20162));
    InMux I__4592 (
            .O(N__20177),
            .I(N__20162));
    InMux I__4591 (
            .O(N__20174),
            .I(N__20162));
    InMux I__4590 (
            .O(N__20173),
            .I(N__20157));
    InMux I__4589 (
            .O(N__20172),
            .I(N__20157));
    Span4Mux_h I__4588 (
            .O(N__20169),
            .I(N__20154));
    LocalMux I__4587 (
            .O(N__20162),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__4586 (
            .O(N__20157),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__4585 (
            .O(N__20154),
            .I(\Lab_UT.di_Mtens_1 ));
    InMux I__4584 (
            .O(N__20147),
            .I(N__20131));
    InMux I__4583 (
            .O(N__20146),
            .I(N__20131));
    InMux I__4582 (
            .O(N__20145),
            .I(N__20131));
    InMux I__4581 (
            .O(N__20144),
            .I(N__20131));
    InMux I__4580 (
            .O(N__20143),
            .I(N__20124));
    InMux I__4579 (
            .O(N__20142),
            .I(N__20124));
    InMux I__4578 (
            .O(N__20141),
            .I(N__20124));
    CascadeMux I__4577 (
            .O(N__20140),
            .I(N__20120));
    LocalMux I__4576 (
            .O(N__20131),
            .I(N__20115));
    LocalMux I__4575 (
            .O(N__20124),
            .I(N__20115));
    CascadeMux I__4574 (
            .O(N__20123),
            .I(N__20112));
    InMux I__4573 (
            .O(N__20120),
            .I(N__20104));
    Span4Mux_h I__4572 (
            .O(N__20115),
            .I(N__20101));
    InMux I__4571 (
            .O(N__20112),
            .I(N__20098));
    InMux I__4570 (
            .O(N__20111),
            .I(N__20093));
    InMux I__4569 (
            .O(N__20110),
            .I(N__20093));
    InMux I__4568 (
            .O(N__20109),
            .I(N__20086));
    InMux I__4567 (
            .O(N__20108),
            .I(N__20086));
    InMux I__4566 (
            .O(N__20107),
            .I(N__20086));
    LocalMux I__4565 (
            .O(N__20104),
            .I(N__20083));
    Span4Mux_v I__4564 (
            .O(N__20101),
            .I(N__20080));
    LocalMux I__4563 (
            .O(N__20098),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4562 (
            .O(N__20093),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4561 (
            .O(N__20086),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv12 I__4560 (
            .O(N__20083),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__4559 (
            .O(N__20080),
            .I(\Lab_UT.di_Mtens_0 ));
    CascadeMux I__4558 (
            .O(N__20069),
            .I(\Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_ ));
    InMux I__4557 (
            .O(N__20066),
            .I(N__20060));
    InMux I__4556 (
            .O(N__20065),
            .I(N__20060));
    LocalMux I__4555 (
            .O(N__20060),
            .I(N__20049));
    InMux I__4554 (
            .O(N__20059),
            .I(N__20046));
    InMux I__4553 (
            .O(N__20058),
            .I(N__20043));
    InMux I__4552 (
            .O(N__20057),
            .I(N__20034));
    InMux I__4551 (
            .O(N__20056),
            .I(N__20034));
    InMux I__4550 (
            .O(N__20055),
            .I(N__20034));
    InMux I__4549 (
            .O(N__20054),
            .I(N__20034));
    InMux I__4548 (
            .O(N__20053),
            .I(N__20025));
    InMux I__4547 (
            .O(N__20052),
            .I(N__20025));
    Span4Mux_v I__4546 (
            .O(N__20049),
            .I(N__20014));
    LocalMux I__4545 (
            .O(N__20046),
            .I(N__20014));
    LocalMux I__4544 (
            .O(N__20043),
            .I(N__20011));
    LocalMux I__4543 (
            .O(N__20034),
            .I(N__20008));
    InMux I__4542 (
            .O(N__20033),
            .I(N__19999));
    InMux I__4541 (
            .O(N__20032),
            .I(N__19999));
    InMux I__4540 (
            .O(N__20031),
            .I(N__19999));
    InMux I__4539 (
            .O(N__20030),
            .I(N__19999));
    LocalMux I__4538 (
            .O(N__20025),
            .I(N__19996));
    InMux I__4537 (
            .O(N__20024),
            .I(N__19989));
    InMux I__4536 (
            .O(N__20023),
            .I(N__19989));
    InMux I__4535 (
            .O(N__20022),
            .I(N__19989));
    InMux I__4534 (
            .O(N__20021),
            .I(N__19982));
    InMux I__4533 (
            .O(N__20020),
            .I(N__19982));
    InMux I__4532 (
            .O(N__20019),
            .I(N__19982));
    Span4Mux_v I__4531 (
            .O(N__20014),
            .I(N__19971));
    Span4Mux_v I__4530 (
            .O(N__20011),
            .I(N__19968));
    Span4Mux_v I__4529 (
            .O(N__20008),
            .I(N__19963));
    LocalMux I__4528 (
            .O(N__19999),
            .I(N__19963));
    Span4Mux_v I__4527 (
            .O(N__19996),
            .I(N__19956));
    LocalMux I__4526 (
            .O(N__19989),
            .I(N__19956));
    LocalMux I__4525 (
            .O(N__19982),
            .I(N__19956));
    InMux I__4524 (
            .O(N__19981),
            .I(N__19953));
    InMux I__4523 (
            .O(N__19980),
            .I(N__19950));
    InMux I__4522 (
            .O(N__19979),
            .I(N__19937));
    InMux I__4521 (
            .O(N__19978),
            .I(N__19937));
    InMux I__4520 (
            .O(N__19977),
            .I(N__19937));
    InMux I__4519 (
            .O(N__19976),
            .I(N__19937));
    InMux I__4518 (
            .O(N__19975),
            .I(N__19937));
    InMux I__4517 (
            .O(N__19974),
            .I(N__19937));
    Odrv4 I__4516 (
            .O(N__19971),
            .I(\Lab_UT.Run ));
    Odrv4 I__4515 (
            .O(N__19968),
            .I(\Lab_UT.Run ));
    Odrv4 I__4514 (
            .O(N__19963),
            .I(\Lab_UT.Run ));
    Odrv4 I__4513 (
            .O(N__19956),
            .I(\Lab_UT.Run ));
    LocalMux I__4512 (
            .O(N__19953),
            .I(\Lab_UT.Run ));
    LocalMux I__4511 (
            .O(N__19950),
            .I(\Lab_UT.Run ));
    LocalMux I__4510 (
            .O(N__19937),
            .I(\Lab_UT.Run ));
    InMux I__4509 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__4508 (
            .O(N__19919),
            .I(N__19916));
    Span4Mux_h I__4507 (
            .O(N__19916),
            .I(N__19913));
    Odrv4 I__4506 (
            .O(N__19913),
            .I(\uu2.bitmapZ0Z_290 ));
    InMux I__4505 (
            .O(N__19910),
            .I(N__19898));
    InMux I__4504 (
            .O(N__19909),
            .I(N__19898));
    InMux I__4503 (
            .O(N__19908),
            .I(N__19898));
    InMux I__4502 (
            .O(N__19907),
            .I(N__19898));
    LocalMux I__4501 (
            .O(N__19898),
            .I(N__19895));
    Odrv4 I__4500 (
            .O(N__19895),
            .I(\Lab_UT.dictrl.N_39_mux ));
    InMux I__4499 (
            .O(N__19892),
            .I(N__19889));
    LocalMux I__4498 (
            .O(N__19889),
            .I(N__19886));
    Span4Mux_h I__4497 (
            .O(N__19886),
            .I(N__19883));
    Odrv4 I__4496 (
            .O(N__19883),
            .I(\Lab_UT.dictrl.g0_0_a3_2 ));
    InMux I__4495 (
            .O(N__19880),
            .I(N__19867));
    CascadeMux I__4494 (
            .O(N__19879),
            .I(N__19864));
    CascadeMux I__4493 (
            .O(N__19878),
            .I(N__19860));
    InMux I__4492 (
            .O(N__19877),
            .I(N__19857));
    InMux I__4491 (
            .O(N__19876),
            .I(N__19852));
    InMux I__4490 (
            .O(N__19875),
            .I(N__19849));
    InMux I__4489 (
            .O(N__19874),
            .I(N__19846));
    InMux I__4488 (
            .O(N__19873),
            .I(N__19843));
    InMux I__4487 (
            .O(N__19872),
            .I(N__19840));
    CascadeMux I__4486 (
            .O(N__19871),
            .I(N__19837));
    CascadeMux I__4485 (
            .O(N__19870),
            .I(N__19834));
    LocalMux I__4484 (
            .O(N__19867),
            .I(N__19829));
    InMux I__4483 (
            .O(N__19864),
            .I(N__19826));
    InMux I__4482 (
            .O(N__19863),
            .I(N__19821));
    InMux I__4481 (
            .O(N__19860),
            .I(N__19821));
    LocalMux I__4480 (
            .O(N__19857),
            .I(N__19818));
    InMux I__4479 (
            .O(N__19856),
            .I(N__19815));
    CascadeMux I__4478 (
            .O(N__19855),
            .I(N__19812));
    LocalMux I__4477 (
            .O(N__19852),
            .I(N__19805));
    LocalMux I__4476 (
            .O(N__19849),
            .I(N__19805));
    LocalMux I__4475 (
            .O(N__19846),
            .I(N__19805));
    LocalMux I__4474 (
            .O(N__19843),
            .I(N__19800));
    LocalMux I__4473 (
            .O(N__19840),
            .I(N__19800));
    InMux I__4472 (
            .O(N__19837),
            .I(N__19797));
    InMux I__4471 (
            .O(N__19834),
            .I(N__19792));
    InMux I__4470 (
            .O(N__19833),
            .I(N__19792));
    InMux I__4469 (
            .O(N__19832),
            .I(N__19789));
    Span4Mux_v I__4468 (
            .O(N__19829),
            .I(N__19784));
    LocalMux I__4467 (
            .O(N__19826),
            .I(N__19784));
    LocalMux I__4466 (
            .O(N__19821),
            .I(N__19781));
    Span4Mux_v I__4465 (
            .O(N__19818),
            .I(N__19775));
    LocalMux I__4464 (
            .O(N__19815),
            .I(N__19772));
    InMux I__4463 (
            .O(N__19812),
            .I(N__19769));
    Span4Mux_v I__4462 (
            .O(N__19805),
            .I(N__19766));
    Span4Mux_h I__4461 (
            .O(N__19800),
            .I(N__19759));
    LocalMux I__4460 (
            .O(N__19797),
            .I(N__19759));
    LocalMux I__4459 (
            .O(N__19792),
            .I(N__19759));
    LocalMux I__4458 (
            .O(N__19789),
            .I(N__19756));
    Span4Mux_h I__4457 (
            .O(N__19784),
            .I(N__19753));
    Span4Mux_v I__4456 (
            .O(N__19781),
            .I(N__19750));
    InMux I__4455 (
            .O(N__19780),
            .I(N__19747));
    InMux I__4454 (
            .O(N__19779),
            .I(N__19742));
    InMux I__4453 (
            .O(N__19778),
            .I(N__19742));
    Span4Mux_h I__4452 (
            .O(N__19775),
            .I(N__19735));
    Span4Mux_h I__4451 (
            .O(N__19772),
            .I(N__19735));
    LocalMux I__4450 (
            .O(N__19769),
            .I(N__19735));
    Span4Mux_h I__4449 (
            .O(N__19766),
            .I(N__19730));
    Span4Mux_v I__4448 (
            .O(N__19759),
            .I(N__19730));
    Span4Mux_s2_v I__4447 (
            .O(N__19756),
            .I(N__19723));
    Span4Mux_v I__4446 (
            .O(N__19753),
            .I(N__19723));
    Span4Mux_h I__4445 (
            .O(N__19750),
            .I(N__19723));
    LocalMux I__4444 (
            .O(N__19747),
            .I(bu_rx_data_2));
    LocalMux I__4443 (
            .O(N__19742),
            .I(bu_rx_data_2));
    Odrv4 I__4442 (
            .O(N__19735),
            .I(bu_rx_data_2));
    Odrv4 I__4441 (
            .O(N__19730),
            .I(bu_rx_data_2));
    Odrv4 I__4440 (
            .O(N__19723),
            .I(bu_rx_data_2));
    CascadeMux I__4439 (
            .O(N__19712),
            .I(N__19709));
    InMux I__4438 (
            .O(N__19709),
            .I(N__19700));
    InMux I__4437 (
            .O(N__19708),
            .I(N__19700));
    InMux I__4436 (
            .O(N__19707),
            .I(N__19700));
    LocalMux I__4435 (
            .O(N__19700),
            .I(N__19695));
    CascadeMux I__4434 (
            .O(N__19699),
            .I(N__19691));
    CascadeMux I__4433 (
            .O(N__19698),
            .I(N__19688));
    Span4Mux_h I__4432 (
            .O(N__19695),
            .I(N__19685));
    InMux I__4431 (
            .O(N__19694),
            .I(N__19678));
    InMux I__4430 (
            .O(N__19691),
            .I(N__19678));
    InMux I__4429 (
            .O(N__19688),
            .I(N__19678));
    Odrv4 I__4428 (
            .O(N__19685),
            .I(bu_rx_data_3_rep1));
    LocalMux I__4427 (
            .O(N__19678),
            .I(bu_rx_data_3_rep1));
    InMux I__4426 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__4425 (
            .O(N__19670),
            .I(N__19667));
    Odrv4 I__4424 (
            .O(N__19667),
            .I(\uu2.bitmapZ0Z_34 ));
    InMux I__4423 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__4422 (
            .O(N__19661),
            .I(N__19658));
    Odrv4 I__4421 (
            .O(N__19658),
            .I(\uu2.bitmapZ0Z_162 ));
    InMux I__4420 (
            .O(N__19655),
            .I(N__19652));
    LocalMux I__4419 (
            .O(N__19652),
            .I(N__19649));
    Odrv4 I__4418 (
            .O(N__19649),
            .I(\Lab_UT.bcd2segment4.segment_0Z0Z_2 ));
    InMux I__4417 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__4416 (
            .O(N__19643),
            .I(N__19640));
    Odrv4 I__4415 (
            .O(N__19640),
            .I(\Lab_UT.bcd2segment4.segmentUQ_0_4 ));
    InMux I__4414 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__4413 (
            .O(N__19634),
            .I(N__19631));
    Odrv4 I__4412 (
            .O(N__19631),
            .I(\Lab_UT.bcd2segment4.segmentUQ_0_5 ));
    InMux I__4411 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__4410 (
            .O(N__19625),
            .I(N__19622));
    Odrv4 I__4409 (
            .O(N__19622),
            .I(\Lab_UT.bcd2segment4.segmentUQ_0_6 ));
    InMux I__4408 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__4407 (
            .O(N__19616),
            .I(\Lab_UT.dictrl.g1_2_3 ));
    InMux I__4406 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__4405 (
            .O(N__19610),
            .I(\Lab_UT.dictrl.g0_1Z0Z_1 ));
    InMux I__4404 (
            .O(N__19607),
            .I(N__19604));
    LocalMux I__4403 (
            .O(N__19604),
            .I(\Lab_UT.dictrl.g0_i_a3_4 ));
    InMux I__4402 (
            .O(N__19601),
            .I(N__19596));
    CascadeMux I__4401 (
            .O(N__19600),
            .I(N__19589));
    CascadeMux I__4400 (
            .O(N__19599),
            .I(N__19585));
    LocalMux I__4399 (
            .O(N__19596),
            .I(N__19582));
    InMux I__4398 (
            .O(N__19595),
            .I(N__19577));
    InMux I__4397 (
            .O(N__19594),
            .I(N__19577));
    InMux I__4396 (
            .O(N__19593),
            .I(N__19572));
    InMux I__4395 (
            .O(N__19592),
            .I(N__19572));
    InMux I__4394 (
            .O(N__19589),
            .I(N__19565));
    InMux I__4393 (
            .O(N__19588),
            .I(N__19565));
    InMux I__4392 (
            .O(N__19585),
            .I(N__19565));
    Odrv4 I__4391 (
            .O(N__19582),
            .I(bu_rx_data_4_rep1));
    LocalMux I__4390 (
            .O(N__19577),
            .I(bu_rx_data_4_rep1));
    LocalMux I__4389 (
            .O(N__19572),
            .I(bu_rx_data_4_rep1));
    LocalMux I__4388 (
            .O(N__19565),
            .I(bu_rx_data_4_rep1));
    InMux I__4387 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__4386 (
            .O(N__19553),
            .I(N__19549));
    InMux I__4385 (
            .O(N__19552),
            .I(N__19546));
    Span4Mux_h I__4384 (
            .O(N__19549),
            .I(N__19537));
    LocalMux I__4383 (
            .O(N__19546),
            .I(N__19534));
    InMux I__4382 (
            .O(N__19545),
            .I(N__19527));
    InMux I__4381 (
            .O(N__19544),
            .I(N__19527));
    InMux I__4380 (
            .O(N__19543),
            .I(N__19527));
    InMux I__4379 (
            .O(N__19542),
            .I(N__19520));
    InMux I__4378 (
            .O(N__19541),
            .I(N__19520));
    InMux I__4377 (
            .O(N__19540),
            .I(N__19520));
    Odrv4 I__4376 (
            .O(N__19537),
            .I(bu_rx_data_7_rep1));
    Odrv12 I__4375 (
            .O(N__19534),
            .I(bu_rx_data_7_rep1));
    LocalMux I__4374 (
            .O(N__19527),
            .I(bu_rx_data_7_rep1));
    LocalMux I__4373 (
            .O(N__19520),
            .I(bu_rx_data_7_rep1));
    InMux I__4372 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__4371 (
            .O(N__19508),
            .I(\Lab_UT.dictrl.g1_4_0 ));
    CascadeMux I__4370 (
            .O(N__19505),
            .I(N__19500));
    InMux I__4369 (
            .O(N__19504),
            .I(N__19496));
    InMux I__4368 (
            .O(N__19503),
            .I(N__19493));
    InMux I__4367 (
            .O(N__19500),
            .I(N__19490));
    CascadeMux I__4366 (
            .O(N__19499),
            .I(N__19487));
    LocalMux I__4365 (
            .O(N__19496),
            .I(N__19481));
    LocalMux I__4364 (
            .O(N__19493),
            .I(N__19481));
    LocalMux I__4363 (
            .O(N__19490),
            .I(N__19478));
    InMux I__4362 (
            .O(N__19487),
            .I(N__19475));
    InMux I__4361 (
            .O(N__19486),
            .I(N__19472));
    Span4Mux_h I__4360 (
            .O(N__19481),
            .I(N__19469));
    Odrv4 I__4359 (
            .O(N__19478),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4358 (
            .O(N__19475),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4357 (
            .O(N__19472),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4356 (
            .O(N__19469),
            .I(bu_rx_data_2_rep1));
    InMux I__4355 (
            .O(N__19460),
            .I(N__19457));
    LocalMux I__4354 (
            .O(N__19457),
            .I(N__19454));
    Span4Mux_h I__4353 (
            .O(N__19454),
            .I(N__19446));
    InMux I__4352 (
            .O(N__19453),
            .I(N__19443));
    InMux I__4351 (
            .O(N__19452),
            .I(N__19438));
    InMux I__4350 (
            .O(N__19451),
            .I(N__19438));
    InMux I__4349 (
            .O(N__19450),
            .I(N__19433));
    InMux I__4348 (
            .O(N__19449),
            .I(N__19433));
    Odrv4 I__4347 (
            .O(N__19446),
            .I(bu_rx_data_fast_2));
    LocalMux I__4346 (
            .O(N__19443),
            .I(bu_rx_data_fast_2));
    LocalMux I__4345 (
            .O(N__19438),
            .I(bu_rx_data_fast_2));
    LocalMux I__4344 (
            .O(N__19433),
            .I(bu_rx_data_fast_2));
    CascadeMux I__4343 (
            .O(N__19424),
            .I(N__19420));
    InMux I__4342 (
            .O(N__19423),
            .I(N__19415));
    InMux I__4341 (
            .O(N__19420),
            .I(N__19408));
    InMux I__4340 (
            .O(N__19419),
            .I(N__19403));
    CascadeMux I__4339 (
            .O(N__19418),
            .I(N__19399));
    LocalMux I__4338 (
            .O(N__19415),
            .I(N__19396));
    InMux I__4337 (
            .O(N__19414),
            .I(N__19393));
    CascadeMux I__4336 (
            .O(N__19413),
            .I(N__19390));
    InMux I__4335 (
            .O(N__19412),
            .I(N__19386));
    InMux I__4334 (
            .O(N__19411),
            .I(N__19383));
    LocalMux I__4333 (
            .O(N__19408),
            .I(N__19380));
    InMux I__4332 (
            .O(N__19407),
            .I(N__19377));
    InMux I__4331 (
            .O(N__19406),
            .I(N__19374));
    LocalMux I__4330 (
            .O(N__19403),
            .I(N__19371));
    InMux I__4329 (
            .O(N__19402),
            .I(N__19366));
    InMux I__4328 (
            .O(N__19399),
            .I(N__19366));
    Span4Mux_v I__4327 (
            .O(N__19396),
            .I(N__19359));
    LocalMux I__4326 (
            .O(N__19393),
            .I(N__19359));
    InMux I__4325 (
            .O(N__19390),
            .I(N__19356));
    InMux I__4324 (
            .O(N__19389),
            .I(N__19353));
    LocalMux I__4323 (
            .O(N__19386),
            .I(N__19347));
    LocalMux I__4322 (
            .O(N__19383),
            .I(N__19347));
    Span4Mux_v I__4321 (
            .O(N__19380),
            .I(N__19340));
    LocalMux I__4320 (
            .O(N__19377),
            .I(N__19340));
    LocalMux I__4319 (
            .O(N__19374),
            .I(N__19340));
    Span4Mux_h I__4318 (
            .O(N__19371),
            .I(N__19333));
    LocalMux I__4317 (
            .O(N__19366),
            .I(N__19333));
    InMux I__4316 (
            .O(N__19365),
            .I(N__19330));
    InMux I__4315 (
            .O(N__19364),
            .I(N__19327));
    Span4Mux_h I__4314 (
            .O(N__19359),
            .I(N__19317));
    LocalMux I__4313 (
            .O(N__19356),
            .I(N__19317));
    LocalMux I__4312 (
            .O(N__19353),
            .I(N__19314));
    InMux I__4311 (
            .O(N__19352),
            .I(N__19311));
    Span4Mux_v I__4310 (
            .O(N__19347),
            .I(N__19306));
    Span4Mux_h I__4309 (
            .O(N__19340),
            .I(N__19306));
    InMux I__4308 (
            .O(N__19339),
            .I(N__19301));
    InMux I__4307 (
            .O(N__19338),
            .I(N__19301));
    Span4Mux_h I__4306 (
            .O(N__19333),
            .I(N__19294));
    LocalMux I__4305 (
            .O(N__19330),
            .I(N__19294));
    LocalMux I__4304 (
            .O(N__19327),
            .I(N__19294));
    InMux I__4303 (
            .O(N__19326),
            .I(N__19291));
    InMux I__4302 (
            .O(N__19325),
            .I(N__19282));
    InMux I__4301 (
            .O(N__19324),
            .I(N__19282));
    InMux I__4300 (
            .O(N__19323),
            .I(N__19282));
    InMux I__4299 (
            .O(N__19322),
            .I(N__19282));
    Span4Mux_v I__4298 (
            .O(N__19317),
            .I(N__19279));
    Sp12to4 I__4297 (
            .O(N__19314),
            .I(N__19270));
    LocalMux I__4296 (
            .O(N__19311),
            .I(N__19270));
    Sp12to4 I__4295 (
            .O(N__19306),
            .I(N__19270));
    LocalMux I__4294 (
            .O(N__19301),
            .I(N__19270));
    Span4Mux_v I__4293 (
            .O(N__19294),
            .I(N__19265));
    LocalMux I__4292 (
            .O(N__19291),
            .I(N__19265));
    LocalMux I__4291 (
            .O(N__19282),
            .I(bu_rx_data_3));
    Odrv4 I__4290 (
            .O(N__19279),
            .I(bu_rx_data_3));
    Odrv12 I__4289 (
            .O(N__19270),
            .I(bu_rx_data_3));
    Odrv4 I__4288 (
            .O(N__19265),
            .I(bu_rx_data_3));
    InMux I__4287 (
            .O(N__19256),
            .I(N__19253));
    LocalMux I__4286 (
            .O(N__19253),
            .I(N__19250));
    Span4Mux_h I__4285 (
            .O(N__19250),
            .I(N__19242));
    InMux I__4284 (
            .O(N__19249),
            .I(N__19239));
    InMux I__4283 (
            .O(N__19248),
            .I(N__19234));
    InMux I__4282 (
            .O(N__19247),
            .I(N__19234));
    InMux I__4281 (
            .O(N__19246),
            .I(N__19229));
    InMux I__4280 (
            .O(N__19245),
            .I(N__19229));
    Odrv4 I__4279 (
            .O(N__19242),
            .I(bu_rx_data_fast_1));
    LocalMux I__4278 (
            .O(N__19239),
            .I(bu_rx_data_fast_1));
    LocalMux I__4277 (
            .O(N__19234),
            .I(bu_rx_data_fast_1));
    LocalMux I__4276 (
            .O(N__19229),
            .I(bu_rx_data_fast_1));
    CascadeMux I__4275 (
            .O(N__19220),
            .I(\Lab_UT.dictrl.g0_i_a3_0_0_cascade_ ));
    CascadeMux I__4274 (
            .O(N__19217),
            .I(\Lab_UT.dictrl.g0_i_a3_0_6_cascade_ ));
    InMux I__4273 (
            .O(N__19214),
            .I(N__19211));
    LocalMux I__4272 (
            .O(N__19211),
            .I(\Lab_UT.dictrl.g0_i_a3_0_5 ));
    InMux I__4271 (
            .O(N__19208),
            .I(N__19202));
    InMux I__4270 (
            .O(N__19207),
            .I(N__19202));
    LocalMux I__4269 (
            .O(N__19202),
            .I(N__19197));
    InMux I__4268 (
            .O(N__19201),
            .I(N__19194));
    InMux I__4267 (
            .O(N__19200),
            .I(N__19191));
    Odrv4 I__4266 (
            .O(N__19197),
            .I(\Lab_UT.dictrl.N_3 ));
    LocalMux I__4265 (
            .O(N__19194),
            .I(\Lab_UT.dictrl.N_3 ));
    LocalMux I__4264 (
            .O(N__19191),
            .I(\Lab_UT.dictrl.N_3 ));
    InMux I__4263 (
            .O(N__19184),
            .I(N__19181));
    LocalMux I__4262 (
            .O(N__19181),
            .I(\Lab_UT.dictrl.g1_4 ));
    CascadeMux I__4261 (
            .O(N__19178),
            .I(N__19172));
    InMux I__4260 (
            .O(N__19177),
            .I(N__19167));
    InMux I__4259 (
            .O(N__19176),
            .I(N__19167));
    InMux I__4258 (
            .O(N__19175),
            .I(N__19164));
    InMux I__4257 (
            .O(N__19172),
            .I(N__19161));
    LocalMux I__4256 (
            .O(N__19167),
            .I(N__19157));
    LocalMux I__4255 (
            .O(N__19164),
            .I(N__19152));
    LocalMux I__4254 (
            .O(N__19161),
            .I(N__19152));
    InMux I__4253 (
            .O(N__19160),
            .I(N__19149));
    Odrv4 I__4252 (
            .O(N__19157),
            .I(\Lab_UT.dictrl.gZ0Z1 ));
    Odrv4 I__4251 (
            .O(N__19152),
            .I(\Lab_UT.dictrl.gZ0Z1 ));
    LocalMux I__4250 (
            .O(N__19149),
            .I(\Lab_UT.dictrl.gZ0Z1 ));
    InMux I__4249 (
            .O(N__19142),
            .I(N__19134));
    InMux I__4248 (
            .O(N__19141),
            .I(N__19131));
    InMux I__4247 (
            .O(N__19140),
            .I(N__19128));
    InMux I__4246 (
            .O(N__19139),
            .I(N__19125));
    InMux I__4245 (
            .O(N__19138),
            .I(N__19120));
    InMux I__4244 (
            .O(N__19137),
            .I(N__19120));
    LocalMux I__4243 (
            .O(N__19134),
            .I(N__19115));
    LocalMux I__4242 (
            .O(N__19131),
            .I(N__19115));
    LocalMux I__4241 (
            .O(N__19128),
            .I(N__19112));
    LocalMux I__4240 (
            .O(N__19125),
            .I(N__19109));
    LocalMux I__4239 (
            .O(N__19120),
            .I(N__19106));
    Span4Mux_v I__4238 (
            .O(N__19115),
            .I(N__19103));
    Odrv4 I__4237 (
            .O(N__19112),
            .I(\Lab_UT.dictrl.next_state12_1 ));
    Odrv4 I__4236 (
            .O(N__19109),
            .I(\Lab_UT.dictrl.next_state12_1 ));
    Odrv12 I__4235 (
            .O(N__19106),
            .I(\Lab_UT.dictrl.next_state12_1 ));
    Odrv4 I__4234 (
            .O(N__19103),
            .I(\Lab_UT.dictrl.next_state12_1 ));
    InMux I__4233 (
            .O(N__19094),
            .I(N__19089));
    InMux I__4232 (
            .O(N__19093),
            .I(N__19086));
    InMux I__4231 (
            .O(N__19092),
            .I(N__19083));
    LocalMux I__4230 (
            .O(N__19089),
            .I(N__19078));
    LocalMux I__4229 (
            .O(N__19086),
            .I(N__19078));
    LocalMux I__4228 (
            .O(N__19083),
            .I(N__19075));
    Span4Mux_v I__4227 (
            .O(N__19078),
            .I(N__19072));
    Odrv4 I__4226 (
            .O(N__19075),
            .I(\Lab_UT.dictrl.next_state32Z0Z_4 ));
    Odrv4 I__4225 (
            .O(N__19072),
            .I(\Lab_UT.dictrl.next_state32Z0Z_4 ));
    CascadeMux I__4224 (
            .O(N__19067),
            .I(\Lab_UT.dictrl.g1Z0Z_0_cascade_ ));
    InMux I__4223 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__4222 (
            .O(N__19061),
            .I(\Lab_UT.dictrl.N_13_0_0 ));
    CascadeMux I__4221 (
            .O(N__19058),
            .I(\Lab_UT.dictrl.g1_2_2_cascade_ ));
    InMux I__4220 (
            .O(N__19055),
            .I(N__19052));
    LocalMux I__4219 (
            .O(N__19052),
            .I(\Lab_UT.dictrl.g2_1_1 ));
    InMux I__4218 (
            .O(N__19049),
            .I(N__19046));
    LocalMux I__4217 (
            .O(N__19046),
            .I(\Lab_UT.dictrl.g2_0 ));
    CascadeMux I__4216 (
            .O(N__19043),
            .I(N__19040));
    InMux I__4215 (
            .O(N__19040),
            .I(N__19037));
    LocalMux I__4214 (
            .O(N__19037),
            .I(N__19033));
    InMux I__4213 (
            .O(N__19036),
            .I(N__19030));
    Odrv4 I__4212 (
            .O(N__19033),
            .I(\Lab_UT.dictrl.i6_mux ));
    LocalMux I__4211 (
            .O(N__19030),
            .I(\Lab_UT.dictrl.i6_mux ));
    CascadeMux I__4210 (
            .O(N__19025),
            .I(\Lab_UT.dictrl.N_15_0_cascade_ ));
    InMux I__4209 (
            .O(N__19022),
            .I(N__19019));
    LocalMux I__4208 (
            .O(N__19019),
            .I(N__19014));
    InMux I__4207 (
            .O(N__19018),
            .I(N__19006));
    InMux I__4206 (
            .O(N__19017),
            .I(N__19006));
    Span4Mux_h I__4205 (
            .O(N__19014),
            .I(N__19002));
    InMux I__4204 (
            .O(N__19013),
            .I(N__18997));
    InMux I__4203 (
            .O(N__19012),
            .I(N__18997));
    InMux I__4202 (
            .O(N__19011),
            .I(N__18994));
    LocalMux I__4201 (
            .O(N__19006),
            .I(N__18991));
    InMux I__4200 (
            .O(N__19005),
            .I(N__18988));
    Odrv4 I__4199 (
            .O(N__19002),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    LocalMux I__4198 (
            .O(N__18997),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    LocalMux I__4197 (
            .O(N__18994),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    Odrv4 I__4196 (
            .O(N__18991),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    LocalMux I__4195 (
            .O(N__18988),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    CascadeMux I__4194 (
            .O(N__18977),
            .I(N__18973));
    CascadeMux I__4193 (
            .O(N__18976),
            .I(N__18970));
    InMux I__4192 (
            .O(N__18973),
            .I(N__18962));
    InMux I__4191 (
            .O(N__18970),
            .I(N__18962));
    InMux I__4190 (
            .O(N__18969),
            .I(N__18955));
    InMux I__4189 (
            .O(N__18968),
            .I(N__18955));
    InMux I__4188 (
            .O(N__18967),
            .I(N__18955));
    LocalMux I__4187 (
            .O(N__18962),
            .I(N__18952));
    LocalMux I__4186 (
            .O(N__18955),
            .I(N__18949));
    Span4Mux_h I__4185 (
            .O(N__18952),
            .I(N__18946));
    Odrv4 I__4184 (
            .O(N__18949),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_0 ));
    Odrv4 I__4183 (
            .O(N__18946),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_0 ));
    CascadeMux I__4182 (
            .O(N__18941),
            .I(N__18935));
    InMux I__4181 (
            .O(N__18940),
            .I(N__18931));
    InMux I__4180 (
            .O(N__18939),
            .I(N__18926));
    InMux I__4179 (
            .O(N__18938),
            .I(N__18926));
    InMux I__4178 (
            .O(N__18935),
            .I(N__18921));
    InMux I__4177 (
            .O(N__18934),
            .I(N__18921));
    LocalMux I__4176 (
            .O(N__18931),
            .I(N__18918));
    LocalMux I__4175 (
            .O(N__18926),
            .I(N__18915));
    LocalMux I__4174 (
            .O(N__18921),
            .I(N__18912));
    Span4Mux_v I__4173 (
            .O(N__18918),
            .I(N__18905));
    Span4Mux_v I__4172 (
            .O(N__18915),
            .I(N__18905));
    Span4Mux_h I__4171 (
            .O(N__18912),
            .I(N__18905));
    Odrv4 I__4170 (
            .O(N__18905),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__4169 (
            .O(N__18902),
            .I(\Lab_UT.dictrl.g0_6_o3_2_0_cascade_ ));
    CascadeMux I__4168 (
            .O(N__18899),
            .I(\Lab_UT.dictrl.N_5_0_cascade_ ));
    InMux I__4167 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__4166 (
            .O(N__18893),
            .I(\Lab_UT.dictrl.g1_3_0 ));
    InMux I__4165 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__4164 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_h I__4163 (
            .O(N__18884),
            .I(N__18881));
    Odrv4 I__4162 (
            .O(N__18881),
            .I(\Lab_UT.dictrl.g2_2 ));
    InMux I__4161 (
            .O(N__18878),
            .I(N__18872));
    InMux I__4160 (
            .O(N__18877),
            .I(N__18867));
    InMux I__4159 (
            .O(N__18876),
            .I(N__18867));
    InMux I__4158 (
            .O(N__18875),
            .I(N__18864));
    LocalMux I__4157 (
            .O(N__18872),
            .I(N__18859));
    LocalMux I__4156 (
            .O(N__18867),
            .I(N__18859));
    LocalMux I__4155 (
            .O(N__18864),
            .I(N__18856));
    Odrv4 I__4154 (
            .O(N__18859),
            .I(\Lab_UT.dictrl.N_16_0_0 ));
    Odrv4 I__4153 (
            .O(N__18856),
            .I(\Lab_UT.dictrl.N_16_0_0 ));
    CascadeMux I__4152 (
            .O(N__18851),
            .I(\Lab_UT.dictrl.N_19_cascade_ ));
    CascadeMux I__4151 (
            .O(N__18848),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ));
    InMux I__4150 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__4149 (
            .O(N__18842),
            .I(\Lab_UT.dictrl.N_19 ));
    InMux I__4148 (
            .O(N__18839),
            .I(N__18835));
    InMux I__4147 (
            .O(N__18838),
            .I(N__18832));
    LocalMux I__4146 (
            .O(N__18835),
            .I(N__18826));
    LocalMux I__4145 (
            .O(N__18832),
            .I(N__18826));
    InMux I__4144 (
            .O(N__18831),
            .I(N__18823));
    Span4Mux_h I__4143 (
            .O(N__18826),
            .I(N__18820));
    LocalMux I__4142 (
            .O(N__18823),
            .I(\Lab_UT.dictrl.N_11_0_0 ));
    Odrv4 I__4141 (
            .O(N__18820),
            .I(\Lab_UT.dictrl.N_11_0_0 ));
    CascadeMux I__4140 (
            .O(N__18815),
            .I(\Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_ ));
    InMux I__4139 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__4138 (
            .O(N__18809),
            .I(\Lab_UT.dictrl.state_ret_5_RNOZ0Z_1 ));
    InMux I__4137 (
            .O(N__18806),
            .I(N__18799));
    InMux I__4136 (
            .O(N__18805),
            .I(N__18799));
    InMux I__4135 (
            .O(N__18804),
            .I(N__18796));
    LocalMux I__4134 (
            .O(N__18799),
            .I(\Lab_UT.dicRun_1 ));
    LocalMux I__4133 (
            .O(N__18796),
            .I(\Lab_UT.dicRun_1 ));
    InMux I__4132 (
            .O(N__18791),
            .I(N__18788));
    LocalMux I__4131 (
            .O(N__18788),
            .I(N__18785));
    Odrv4 I__4130 (
            .O(N__18785),
            .I(\Lab_UT.dictrl.N_10 ));
    InMux I__4129 (
            .O(N__18782),
            .I(N__18779));
    LocalMux I__4128 (
            .O(N__18779),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_2 ));
    CascadeMux I__4127 (
            .O(N__18776),
            .I(\Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_ ));
    InMux I__4126 (
            .O(N__18773),
            .I(N__18766));
    InMux I__4125 (
            .O(N__18772),
            .I(N__18763));
    InMux I__4124 (
            .O(N__18771),
            .I(N__18760));
    InMux I__4123 (
            .O(N__18770),
            .I(N__18757));
    InMux I__4122 (
            .O(N__18769),
            .I(N__18754));
    LocalMux I__4121 (
            .O(N__18766),
            .I(\Lab_UT.dictrl.N_5 ));
    LocalMux I__4120 (
            .O(N__18763),
            .I(\Lab_UT.dictrl.N_5 ));
    LocalMux I__4119 (
            .O(N__18760),
            .I(\Lab_UT.dictrl.N_5 ));
    LocalMux I__4118 (
            .O(N__18757),
            .I(\Lab_UT.dictrl.N_5 ));
    LocalMux I__4117 (
            .O(N__18754),
            .I(\Lab_UT.dictrl.N_5 ));
    InMux I__4116 (
            .O(N__18743),
            .I(N__18740));
    LocalMux I__4115 (
            .O(N__18740),
            .I(N__18737));
    Odrv4 I__4114 (
            .O(N__18737),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_3 ));
    CascadeMux I__4113 (
            .O(N__18734),
            .I(\Lab_UT.dictrl.N_14_cascade_ ));
    InMux I__4112 (
            .O(N__18731),
            .I(N__18728));
    LocalMux I__4111 (
            .O(N__18728),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_3 ));
    CascadeMux I__4110 (
            .O(N__18725),
            .I(\Lab_UT.dictrl.N_7_cascade_ ));
    CascadeMux I__4109 (
            .O(N__18722),
            .I(\Lab_UT.dictrl.N_13_0_cascade_ ));
    CascadeMux I__4108 (
            .O(N__18719),
            .I(\Lab_UT.dictrl.N_6_cascade_ ));
    CascadeMux I__4107 (
            .O(N__18716),
            .I(N__18713));
    InMux I__4106 (
            .O(N__18713),
            .I(N__18709));
    InMux I__4105 (
            .O(N__18712),
            .I(N__18706));
    LocalMux I__4104 (
            .O(N__18709),
            .I(N__18701));
    LocalMux I__4103 (
            .O(N__18706),
            .I(N__18698));
    CascadeMux I__4102 (
            .O(N__18705),
            .I(N__18695));
    InMux I__4101 (
            .O(N__18704),
            .I(N__18692));
    Span4Mux_v I__4100 (
            .O(N__18701),
            .I(N__18687));
    Span4Mux_s3_v I__4099 (
            .O(N__18698),
            .I(N__18687));
    InMux I__4098 (
            .O(N__18695),
            .I(N__18684));
    LocalMux I__4097 (
            .O(N__18692),
            .I(N__18681));
    Span4Mux_v I__4096 (
            .O(N__18687),
            .I(N__18676));
    LocalMux I__4095 (
            .O(N__18684),
            .I(N__18676));
    Odrv12 I__4094 (
            .O(N__18681),
            .I(\Lab_UT.LdStens ));
    Odrv4 I__4093 (
            .O(N__18676),
            .I(\Lab_UT.LdStens ));
    InMux I__4092 (
            .O(N__18671),
            .I(N__18666));
    InMux I__4091 (
            .O(N__18670),
            .I(N__18661));
    InMux I__4090 (
            .O(N__18669),
            .I(N__18661));
    LocalMux I__4089 (
            .O(N__18666),
            .I(\Lab_UT.state_i_3_2 ));
    LocalMux I__4088 (
            .O(N__18661),
            .I(\Lab_UT.state_i_3_2 ));
    CascadeMux I__4087 (
            .O(N__18656),
            .I(N__18653));
    InMux I__4086 (
            .O(N__18653),
            .I(N__18650));
    LocalMux I__4085 (
            .O(N__18650),
            .I(\Lab_UT.LdStens_i_3 ));
    InMux I__4084 (
            .O(N__18647),
            .I(N__18641));
    InMux I__4083 (
            .O(N__18646),
            .I(N__18641));
    LocalMux I__4082 (
            .O(N__18641),
            .I(N__18638));
    Span4Mux_v I__4081 (
            .O(N__18638),
            .I(N__18635));
    Odrv4 I__4080 (
            .O(N__18635),
            .I(\Lab_UT.didp.ce_10_0_1 ));
    InMux I__4079 (
            .O(N__18632),
            .I(N__18629));
    LocalMux I__4078 (
            .O(N__18629),
            .I(N__18626));
    Span4Mux_v I__4077 (
            .O(N__18626),
            .I(N__18623));
    Span4Mux_h I__4076 (
            .O(N__18623),
            .I(N__18620));
    Odrv4 I__4075 (
            .O(N__18620),
            .I(\Lab_UT.dictrl.m27_1 ));
    InMux I__4074 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__4073 (
            .O(N__18614),
            .I(N__18611));
    Odrv12 I__4072 (
            .O(N__18611),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_0 ));
    InMux I__4071 (
            .O(N__18608),
            .I(N__18605));
    LocalMux I__4070 (
            .O(N__18605),
            .I(N__18602));
    Odrv4 I__4069 (
            .O(N__18602),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_3 ));
    InMux I__4068 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__4067 (
            .O(N__18596),
            .I(N__18593));
    Span4Mux_v I__4066 (
            .O(N__18593),
            .I(N__18590));
    Odrv4 I__4065 (
            .O(N__18590),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_2 ));
    InMux I__4064 (
            .O(N__18587),
            .I(N__18584));
    LocalMux I__4063 (
            .O(N__18584),
            .I(N__18581));
    Odrv4 I__4062 (
            .O(N__18581),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_5 ));
    InMux I__4061 (
            .O(N__18578),
            .I(N__18575));
    LocalMux I__4060 (
            .O(N__18575),
            .I(N__18572));
    Span4Mux_v I__4059 (
            .O(N__18572),
            .I(N__18569));
    Odrv4 I__4058 (
            .O(N__18569),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_6 ));
    InMux I__4057 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__4056 (
            .O(N__18563),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_0 ));
    InMux I__4055 (
            .O(N__18560),
            .I(N__18557));
    LocalMux I__4054 (
            .O(N__18557),
            .I(N__18554));
    Span4Mux_h I__4053 (
            .O(N__18554),
            .I(N__18551));
    Odrv4 I__4052 (
            .O(N__18551),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_1 ));
    InMux I__4051 (
            .O(N__18548),
            .I(N__18527));
    InMux I__4050 (
            .O(N__18547),
            .I(N__18527));
    InMux I__4049 (
            .O(N__18546),
            .I(N__18527));
    InMux I__4048 (
            .O(N__18545),
            .I(N__18527));
    InMux I__4047 (
            .O(N__18544),
            .I(N__18527));
    InMux I__4046 (
            .O(N__18543),
            .I(N__18527));
    InMux I__4045 (
            .O(N__18542),
            .I(N__18527));
    LocalMux I__4044 (
            .O(N__18527),
            .I(N__18520));
    InMux I__4043 (
            .O(N__18526),
            .I(N__18517));
    InMux I__4042 (
            .O(N__18525),
            .I(N__18512));
    InMux I__4041 (
            .O(N__18524),
            .I(N__18512));
    InMux I__4040 (
            .O(N__18523),
            .I(N__18509));
    Span4Mux_h I__4039 (
            .O(N__18520),
            .I(N__18506));
    LocalMux I__4038 (
            .O(N__18517),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__4037 (
            .O(N__18512),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__4036 (
            .O(N__18509),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__4035 (
            .O(N__18506),
            .I(\Lab_UT.di_Sones_2 ));
    CascadeMux I__4034 (
            .O(N__18497),
            .I(N__18491));
    CascadeMux I__4033 (
            .O(N__18496),
            .I(N__18488));
    CascadeMux I__4032 (
            .O(N__18495),
            .I(N__18484));
    InMux I__4031 (
            .O(N__18494),
            .I(N__18466));
    InMux I__4030 (
            .O(N__18491),
            .I(N__18466));
    InMux I__4029 (
            .O(N__18488),
            .I(N__18466));
    InMux I__4028 (
            .O(N__18487),
            .I(N__18466));
    InMux I__4027 (
            .O(N__18484),
            .I(N__18466));
    InMux I__4026 (
            .O(N__18483),
            .I(N__18466));
    InMux I__4025 (
            .O(N__18482),
            .I(N__18466));
    InMux I__4024 (
            .O(N__18481),
            .I(N__18459));
    LocalMux I__4023 (
            .O(N__18466),
            .I(N__18456));
    InMux I__4022 (
            .O(N__18465),
            .I(N__18453));
    InMux I__4021 (
            .O(N__18464),
            .I(N__18448));
    InMux I__4020 (
            .O(N__18463),
            .I(N__18448));
    InMux I__4019 (
            .O(N__18462),
            .I(N__18445));
    LocalMux I__4018 (
            .O(N__18459),
            .I(N__18440));
    Span4Mux_v I__4017 (
            .O(N__18456),
            .I(N__18440));
    LocalMux I__4016 (
            .O(N__18453),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__4015 (
            .O(N__18448),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__4014 (
            .O(N__18445),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__4013 (
            .O(N__18440),
            .I(\Lab_UT.di_Sones_1 ));
    CascadeMux I__4012 (
            .O(N__18431),
            .I(N__18425));
    CascadeMux I__4011 (
            .O(N__18430),
            .I(N__18422));
    CascadeMux I__4010 (
            .O(N__18429),
            .I(N__18419));
    CascadeMux I__4009 (
            .O(N__18428),
            .I(N__18416));
    InMux I__4008 (
            .O(N__18425),
            .I(N__18398));
    InMux I__4007 (
            .O(N__18422),
            .I(N__18398));
    InMux I__4006 (
            .O(N__18419),
            .I(N__18398));
    InMux I__4005 (
            .O(N__18416),
            .I(N__18398));
    InMux I__4004 (
            .O(N__18415),
            .I(N__18398));
    InMux I__4003 (
            .O(N__18414),
            .I(N__18398));
    InMux I__4002 (
            .O(N__18413),
            .I(N__18398));
    LocalMux I__4001 (
            .O(N__18398),
            .I(N__18392));
    InMux I__4000 (
            .O(N__18397),
            .I(N__18389));
    InMux I__3999 (
            .O(N__18396),
            .I(N__18386));
    InMux I__3998 (
            .O(N__18395),
            .I(N__18383));
    Span4Mux_h I__3997 (
            .O(N__18392),
            .I(N__18380));
    LocalMux I__3996 (
            .O(N__18389),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3995 (
            .O(N__18386),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3994 (
            .O(N__18383),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv4 I__3993 (
            .O(N__18380),
            .I(\Lab_UT.di_Sones_3 ));
    InMux I__3992 (
            .O(N__18371),
            .I(N__18349));
    InMux I__3991 (
            .O(N__18370),
            .I(N__18349));
    InMux I__3990 (
            .O(N__18369),
            .I(N__18349));
    InMux I__3989 (
            .O(N__18368),
            .I(N__18349));
    InMux I__3988 (
            .O(N__18367),
            .I(N__18349));
    InMux I__3987 (
            .O(N__18366),
            .I(N__18349));
    InMux I__3986 (
            .O(N__18365),
            .I(N__18349));
    CascadeMux I__3985 (
            .O(N__18364),
            .I(N__18341));
    LocalMux I__3984 (
            .O(N__18349),
            .I(N__18338));
    InMux I__3983 (
            .O(N__18348),
            .I(N__18331));
    InMux I__3982 (
            .O(N__18347),
            .I(N__18331));
    InMux I__3981 (
            .O(N__18346),
            .I(N__18331));
    InMux I__3980 (
            .O(N__18345),
            .I(N__18328));
    InMux I__3979 (
            .O(N__18344),
            .I(N__18323));
    InMux I__3978 (
            .O(N__18341),
            .I(N__18323));
    Span4Mux_h I__3977 (
            .O(N__18338),
            .I(N__18320));
    LocalMux I__3976 (
            .O(N__18331),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3975 (
            .O(N__18328),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3974 (
            .O(N__18323),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__3973 (
            .O(N__18320),
            .I(\Lab_UT.di_Sones_0 ));
    CascadeMux I__3972 (
            .O(N__18311),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ));
    InMux I__3971 (
            .O(N__18308),
            .I(N__18305));
    LocalMux I__3970 (
            .O(N__18305),
            .I(N__18302));
    Odrv4 I__3969 (
            .O(N__18302),
            .I(\uu2.bitmapZ0Z_218 ));
    CascadeMux I__3968 (
            .O(N__18299),
            .I(\uu2.mem0.bitmap_pmux_16_ns_1_cascade_ ));
    InMux I__3967 (
            .O(N__18296),
            .I(N__18293));
    LocalMux I__3966 (
            .O(N__18293),
            .I(N__18289));
    InMux I__3965 (
            .O(N__18292),
            .I(N__18285));
    Span4Mux_h I__3964 (
            .O(N__18289),
            .I(N__18281));
    InMux I__3963 (
            .O(N__18288),
            .I(N__18278));
    LocalMux I__3962 (
            .O(N__18285),
            .I(N__18275));
    InMux I__3961 (
            .O(N__18284),
            .I(N__18272));
    Odrv4 I__3960 (
            .O(N__18281),
            .I(\uu2.N_30_i ));
    LocalMux I__3959 (
            .O(N__18278),
            .I(\uu2.N_30_i ));
    Odrv12 I__3958 (
            .O(N__18275),
            .I(\uu2.N_30_i ));
    LocalMux I__3957 (
            .O(N__18272),
            .I(\uu2.N_30_i ));
    CascadeMux I__3956 (
            .O(N__18263),
            .I(\uu2.mem0.N_22_cascade_ ));
    InMux I__3955 (
            .O(N__18260),
            .I(N__18257));
    LocalMux I__3954 (
            .O(N__18257),
            .I(N__18254));
    Odrv4 I__3953 (
            .O(N__18254),
            .I(\uu2.mem0.G_11_0_0_a3_6_0 ));
    InMux I__3952 (
            .O(N__18251),
            .I(N__18245));
    InMux I__3951 (
            .O(N__18250),
            .I(N__18245));
    LocalMux I__3950 (
            .O(N__18245),
            .I(\uu2.bitmapZ0Z_200 ));
    CascadeMux I__3949 (
            .O(N__18242),
            .I(N__18238));
    InMux I__3948 (
            .O(N__18241),
            .I(N__18232));
    InMux I__3947 (
            .O(N__18238),
            .I(N__18227));
    InMux I__3946 (
            .O(N__18237),
            .I(N__18227));
    CascadeMux I__3945 (
            .O(N__18236),
            .I(N__18223));
    InMux I__3944 (
            .O(N__18235),
            .I(N__18220));
    LocalMux I__3943 (
            .O(N__18232),
            .I(N__18215));
    LocalMux I__3942 (
            .O(N__18227),
            .I(N__18215));
    InMux I__3941 (
            .O(N__18226),
            .I(N__18212));
    InMux I__3940 (
            .O(N__18223),
            .I(N__18209));
    LocalMux I__3939 (
            .O(N__18220),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__3938 (
            .O(N__18215),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__3937 (
            .O(N__18212),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__3936 (
            .O(N__18209),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    CascadeMux I__3935 (
            .O(N__18200),
            .I(N__18197));
    InMux I__3934 (
            .O(N__18197),
            .I(N__18191));
    InMux I__3933 (
            .O(N__18196),
            .I(N__18191));
    LocalMux I__3932 (
            .O(N__18191),
            .I(\uu2.bitmapZ0Z_72 ));
    CascadeMux I__3931 (
            .O(N__18188),
            .I(N__18184));
    InMux I__3930 (
            .O(N__18187),
            .I(N__18176));
    InMux I__3929 (
            .O(N__18184),
            .I(N__18173));
    InMux I__3928 (
            .O(N__18183),
            .I(N__18170));
    InMux I__3927 (
            .O(N__18182),
            .I(N__18165));
    InMux I__3926 (
            .O(N__18181),
            .I(N__18165));
    InMux I__3925 (
            .O(N__18180),
            .I(N__18160));
    InMux I__3924 (
            .O(N__18179),
            .I(N__18160));
    LocalMux I__3923 (
            .O(N__18176),
            .I(N__18157));
    LocalMux I__3922 (
            .O(N__18173),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3921 (
            .O(N__18170),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3920 (
            .O(N__18165),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3919 (
            .O(N__18160),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__3918 (
            .O(N__18157),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    InMux I__3917 (
            .O(N__18146),
            .I(N__18140));
    InMux I__3916 (
            .O(N__18145),
            .I(N__18140));
    LocalMux I__3915 (
            .O(N__18140),
            .I(N__18137));
    Odrv4 I__3914 (
            .O(N__18137),
            .I(\uu2.bitmapZ0Z_203 ));
    CascadeMux I__3913 (
            .O(N__18134),
            .I(\uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_ ));
    InMux I__3912 (
            .O(N__18131),
            .I(N__18127));
    InMux I__3911 (
            .O(N__18130),
            .I(N__18124));
    LocalMux I__3910 (
            .O(N__18127),
            .I(\uu2.bitmapZ0Z_75 ));
    LocalMux I__3909 (
            .O(N__18124),
            .I(\uu2.bitmapZ0Z_75 ));
    CascadeMux I__3908 (
            .O(N__18119),
            .I(N__18108));
    CascadeMux I__3907 (
            .O(N__18118),
            .I(N__18105));
    CascadeMux I__3906 (
            .O(N__18117),
            .I(N__18099));
    CascadeMux I__3905 (
            .O(N__18116),
            .I(N__18096));
    InMux I__3904 (
            .O(N__18115),
            .I(N__18091));
    InMux I__3903 (
            .O(N__18114),
            .I(N__18091));
    InMux I__3902 (
            .O(N__18113),
            .I(N__18088));
    InMux I__3901 (
            .O(N__18112),
            .I(N__18081));
    InMux I__3900 (
            .O(N__18111),
            .I(N__18081));
    InMux I__3899 (
            .O(N__18108),
            .I(N__18081));
    InMux I__3898 (
            .O(N__18105),
            .I(N__18076));
    InMux I__3897 (
            .O(N__18104),
            .I(N__18076));
    CascadeMux I__3896 (
            .O(N__18103),
            .I(N__18073));
    InMux I__3895 (
            .O(N__18102),
            .I(N__18069));
    InMux I__3894 (
            .O(N__18099),
            .I(N__18066));
    InMux I__3893 (
            .O(N__18096),
            .I(N__18063));
    LocalMux I__3892 (
            .O(N__18091),
            .I(N__18060));
    LocalMux I__3891 (
            .O(N__18088),
            .I(N__18053));
    LocalMux I__3890 (
            .O(N__18081),
            .I(N__18053));
    LocalMux I__3889 (
            .O(N__18076),
            .I(N__18053));
    InMux I__3888 (
            .O(N__18073),
            .I(N__18050));
    InMux I__3887 (
            .O(N__18072),
            .I(N__18047));
    LocalMux I__3886 (
            .O(N__18069),
            .I(N__18042));
    LocalMux I__3885 (
            .O(N__18066),
            .I(N__18042));
    LocalMux I__3884 (
            .O(N__18063),
            .I(N__18033));
    Span4Mux_v I__3883 (
            .O(N__18060),
            .I(N__18033));
    Span4Mux_v I__3882 (
            .O(N__18053),
            .I(N__18033));
    LocalMux I__3881 (
            .O(N__18050),
            .I(N__18033));
    LocalMux I__3880 (
            .O(N__18047),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__3879 (
            .O(N__18042),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__3878 (
            .O(N__18033),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__3877 (
            .O(N__18026),
            .I(N__18022));
    InMux I__3876 (
            .O(N__18025),
            .I(N__18019));
    LocalMux I__3875 (
            .O(N__18022),
            .I(N__18016));
    LocalMux I__3874 (
            .O(N__18019),
            .I(\uu2.N_30_i_1 ));
    Odrv4 I__3873 (
            .O(N__18016),
            .I(\uu2.N_30_i_1 ));
    CascadeMux I__3872 (
            .O(N__18011),
            .I(\uu2.mem0.N_22_0_cascade_ ));
    InMux I__3871 (
            .O(N__18008),
            .I(N__18005));
    LocalMux I__3870 (
            .O(N__18005),
            .I(N__18002));
    Odrv12 I__3869 (
            .O(N__18002),
            .I(\uu2.N_104 ));
    InMux I__3868 (
            .O(N__17999),
            .I(N__17996));
    LocalMux I__3867 (
            .O(N__17996),
            .I(\uu2.mem0.bitmap_pmux_27_ns_1_0 ));
    InMux I__3866 (
            .O(N__17993),
            .I(N__17978));
    InMux I__3865 (
            .O(N__17992),
            .I(N__17978));
    InMux I__3864 (
            .O(N__17991),
            .I(N__17978));
    InMux I__3863 (
            .O(N__17990),
            .I(N__17973));
    InMux I__3862 (
            .O(N__17989),
            .I(N__17970));
    InMux I__3861 (
            .O(N__17988),
            .I(N__17963));
    InMux I__3860 (
            .O(N__17987),
            .I(N__17963));
    InMux I__3859 (
            .O(N__17986),
            .I(N__17963));
    InMux I__3858 (
            .O(N__17985),
            .I(N__17960));
    LocalMux I__3857 (
            .O(N__17978),
            .I(N__17957));
    InMux I__3856 (
            .O(N__17977),
            .I(N__17952));
    InMux I__3855 (
            .O(N__17976),
            .I(N__17952));
    LocalMux I__3854 (
            .O(N__17973),
            .I(N__17947));
    LocalMux I__3853 (
            .O(N__17970),
            .I(N__17947));
    LocalMux I__3852 (
            .O(N__17963),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3851 (
            .O(N__17960),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3850 (
            .O(N__17957),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3849 (
            .O(N__17952),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3848 (
            .O(N__17947),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__3847 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__3846 (
            .O(N__17933),
            .I(\uu2.mem0.N_109 ));
    InMux I__3845 (
            .O(N__17930),
            .I(N__17924));
    InMux I__3844 (
            .O(N__17929),
            .I(N__17924));
    LocalMux I__3843 (
            .O(N__17924),
            .I(\uu2.bitmap_pmux_19_ns_1 ));
    CascadeMux I__3842 (
            .O(N__17921),
            .I(N__17914));
    InMux I__3841 (
            .O(N__17920),
            .I(N__17905));
    InMux I__3840 (
            .O(N__17919),
            .I(N__17905));
    InMux I__3839 (
            .O(N__17918),
            .I(N__17900));
    InMux I__3838 (
            .O(N__17917),
            .I(N__17891));
    InMux I__3837 (
            .O(N__17914),
            .I(N__17891));
    InMux I__3836 (
            .O(N__17913),
            .I(N__17891));
    InMux I__3835 (
            .O(N__17912),
            .I(N__17891));
    CascadeMux I__3834 (
            .O(N__17911),
            .I(N__17885));
    CascadeMux I__3833 (
            .O(N__17910),
            .I(N__17881));
    LocalMux I__3832 (
            .O(N__17905),
            .I(N__17877));
    CascadeMux I__3831 (
            .O(N__17904),
            .I(N__17874));
    InMux I__3830 (
            .O(N__17903),
            .I(N__17871));
    LocalMux I__3829 (
            .O(N__17900),
            .I(N__17866));
    LocalMux I__3828 (
            .O(N__17891),
            .I(N__17866));
    CascadeMux I__3827 (
            .O(N__17890),
            .I(N__17861));
    CascadeMux I__3826 (
            .O(N__17889),
            .I(N__17858));
    InMux I__3825 (
            .O(N__17888),
            .I(N__17855));
    InMux I__3824 (
            .O(N__17885),
            .I(N__17848));
    InMux I__3823 (
            .O(N__17884),
            .I(N__17848));
    InMux I__3822 (
            .O(N__17881),
            .I(N__17848));
    InMux I__3821 (
            .O(N__17880),
            .I(N__17845));
    Span4Mux_v I__3820 (
            .O(N__17877),
            .I(N__17842));
    InMux I__3819 (
            .O(N__17874),
            .I(N__17839));
    LocalMux I__3818 (
            .O(N__17871),
            .I(N__17836));
    Span4Mux_h I__3817 (
            .O(N__17866),
            .I(N__17833));
    InMux I__3816 (
            .O(N__17865),
            .I(N__17824));
    InMux I__3815 (
            .O(N__17864),
            .I(N__17824));
    InMux I__3814 (
            .O(N__17861),
            .I(N__17824));
    InMux I__3813 (
            .O(N__17858),
            .I(N__17824));
    LocalMux I__3812 (
            .O(N__17855),
            .I(N__17821));
    LocalMux I__3811 (
            .O(N__17848),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3810 (
            .O(N__17845),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3809 (
            .O(N__17842),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3808 (
            .O(N__17839),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv12 I__3807 (
            .O(N__17836),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3806 (
            .O(N__17833),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3805 (
            .O(N__17824),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3804 (
            .O(N__17821),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    CascadeMux I__3803 (
            .O(N__17804),
            .I(N__17801));
    InMux I__3802 (
            .O(N__17801),
            .I(N__17795));
    InMux I__3801 (
            .O(N__17800),
            .I(N__17795));
    LocalMux I__3800 (
            .O(N__17795),
            .I(N__17792));
    Span4Mux_s3_h I__3799 (
            .O(N__17792),
            .I(N__17789));
    Odrv4 I__3798 (
            .O(N__17789),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__3797 (
            .O(N__17786),
            .I(N__17782));
    InMux I__3796 (
            .O(N__17785),
            .I(N__17777));
    InMux I__3795 (
            .O(N__17782),
            .I(N__17777));
    LocalMux I__3794 (
            .O(N__17777),
            .I(N__17774));
    Odrv4 I__3793 (
            .O(N__17774),
            .I(\uu2.bitmapZ0Z_93 ));
    InMux I__3792 (
            .O(N__17771),
            .I(N__17768));
    LocalMux I__3791 (
            .O(N__17768),
            .I(\uu2.mem0.N_109_0 ));
    InMux I__3790 (
            .O(N__17765),
            .I(N__17759));
    CascadeMux I__3789 (
            .O(N__17764),
            .I(N__17754));
    CascadeMux I__3788 (
            .O(N__17763),
            .I(N__17751));
    InMux I__3787 (
            .O(N__17762),
            .I(N__17745));
    LocalMux I__3786 (
            .O(N__17759),
            .I(N__17742));
    InMux I__3785 (
            .O(N__17758),
            .I(N__17738));
    InMux I__3784 (
            .O(N__17757),
            .I(N__17735));
    InMux I__3783 (
            .O(N__17754),
            .I(N__17728));
    InMux I__3782 (
            .O(N__17751),
            .I(N__17728));
    InMux I__3781 (
            .O(N__17750),
            .I(N__17728));
    InMux I__3780 (
            .O(N__17749),
            .I(N__17723));
    InMux I__3779 (
            .O(N__17748),
            .I(N__17723));
    LocalMux I__3778 (
            .O(N__17745),
            .I(N__17718));
    Span4Mux_v I__3777 (
            .O(N__17742),
            .I(N__17718));
    InMux I__3776 (
            .O(N__17741),
            .I(N__17715));
    LocalMux I__3775 (
            .O(N__17738),
            .I(N__17710));
    LocalMux I__3774 (
            .O(N__17735),
            .I(N__17710));
    LocalMux I__3773 (
            .O(N__17728),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__3772 (
            .O(N__17723),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv4 I__3771 (
            .O(N__17718),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__3770 (
            .O(N__17715),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv4 I__3769 (
            .O(N__17710),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    CascadeMux I__3768 (
            .O(N__17699),
            .I(N__17696));
    InMux I__3767 (
            .O(N__17696),
            .I(N__17693));
    LocalMux I__3766 (
            .O(N__17693),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__3765 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__3764 (
            .O(N__17687),
            .I(\uu2.bitmapZ0Z_194 ));
    CascadeMux I__3763 (
            .O(N__17684),
            .I(\uu2.bitmap_pmux_20_ns_1_cascade_ ));
    InMux I__3762 (
            .O(N__17681),
            .I(N__17678));
    LocalMux I__3761 (
            .O(N__17678),
            .I(N__17675));
    Odrv4 I__3760 (
            .O(N__17675),
            .I(\uu2.mem0.N_108 ));
    InMux I__3759 (
            .O(N__17672),
            .I(N__17666));
    InMux I__3758 (
            .O(N__17671),
            .I(N__17666));
    LocalMux I__3757 (
            .O(N__17666),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__3756 (
            .O(N__17663),
            .I(N__17657));
    InMux I__3755 (
            .O(N__17662),
            .I(N__17657));
    LocalMux I__3754 (
            .O(N__17657),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__3753 (
            .O(N__17654),
            .I(N__17651));
    LocalMux I__3752 (
            .O(N__17651),
            .I(\uu2.bitmap_pmux_20_ns_1 ));
    CascadeMux I__3751 (
            .O(N__17648),
            .I(\uu2.mem0.N_108_0_cascade_ ));
    InMux I__3750 (
            .O(N__17645),
            .I(N__17642));
    LocalMux I__3749 (
            .O(N__17642),
            .I(N__17639));
    Span4Mux_h I__3748 (
            .O(N__17639),
            .I(N__17636));
    Odrv4 I__3747 (
            .O(N__17636),
            .I(\uu2.mem0.N_404_0 ));
    CascadeMux I__3746 (
            .O(N__17633),
            .I(N__17624));
    InMux I__3745 (
            .O(N__17632),
            .I(N__17619));
    InMux I__3744 (
            .O(N__17631),
            .I(N__17619));
    CascadeMux I__3743 (
            .O(N__17630),
            .I(N__17616));
    InMux I__3742 (
            .O(N__17629),
            .I(N__17612));
    InMux I__3741 (
            .O(N__17628),
            .I(N__17609));
    InMux I__3740 (
            .O(N__17627),
            .I(N__17606));
    InMux I__3739 (
            .O(N__17624),
            .I(N__17603));
    LocalMux I__3738 (
            .O(N__17619),
            .I(N__17600));
    InMux I__3737 (
            .O(N__17616),
            .I(N__17597));
    InMux I__3736 (
            .O(N__17615),
            .I(N__17594));
    LocalMux I__3735 (
            .O(N__17612),
            .I(N__17591));
    LocalMux I__3734 (
            .O(N__17609),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3733 (
            .O(N__17606),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3732 (
            .O(N__17603),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__3731 (
            .O(N__17600),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3730 (
            .O(N__17597),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3729 (
            .O(N__17594),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__3728 (
            .O(N__17591),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    CascadeMux I__3727 (
            .O(N__17576),
            .I(\uu2.N_104_cascade_ ));
    CascadeMux I__3726 (
            .O(N__17573),
            .I(\uu2.mem0.G_11_0_0_a3_5_0_cascade_ ));
    InMux I__3725 (
            .O(N__17570),
            .I(N__17567));
    LocalMux I__3724 (
            .O(N__17567),
            .I(\uu2.mem0.N_40 ));
    InMux I__3723 (
            .O(N__17564),
            .I(N__17561));
    LocalMux I__3722 (
            .O(N__17561),
            .I(\uu2.mem0.N_30 ));
    InMux I__3721 (
            .O(N__17558),
            .I(N__17552));
    InMux I__3720 (
            .O(N__17557),
            .I(N__17552));
    LocalMux I__3719 (
            .O(N__17552),
            .I(N__17548));
    InMux I__3718 (
            .O(N__17551),
            .I(N__17542));
    Span4Mux_h I__3717 (
            .O(N__17548),
            .I(N__17538));
    InMux I__3716 (
            .O(N__17547),
            .I(N__17531));
    InMux I__3715 (
            .O(N__17546),
            .I(N__17531));
    InMux I__3714 (
            .O(N__17545),
            .I(N__17531));
    LocalMux I__3713 (
            .O(N__17542),
            .I(N__17528));
    InMux I__3712 (
            .O(N__17541),
            .I(N__17525));
    Odrv4 I__3711 (
            .O(N__17538),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__3710 (
            .O(N__17531),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__3709 (
            .O(N__17528),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__3708 (
            .O(N__17525),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    InMux I__3707 (
            .O(N__17516),
            .I(N__17508));
    InMux I__3706 (
            .O(N__17515),
            .I(N__17508));
    InMux I__3705 (
            .O(N__17514),
            .I(N__17501));
    InMux I__3704 (
            .O(N__17513),
            .I(N__17501));
    LocalMux I__3703 (
            .O(N__17508),
            .I(N__17498));
    InMux I__3702 (
            .O(N__17507),
            .I(N__17493));
    InMux I__3701 (
            .O(N__17506),
            .I(N__17493));
    LocalMux I__3700 (
            .O(N__17501),
            .I(N__17477));
    Span4Mux_v I__3699 (
            .O(N__17498),
            .I(N__17477));
    LocalMux I__3698 (
            .O(N__17493),
            .I(N__17477));
    InMux I__3697 (
            .O(N__17492),
            .I(N__17473));
    InMux I__3696 (
            .O(N__17491),
            .I(N__17468));
    InMux I__3695 (
            .O(N__17490),
            .I(N__17468));
    InMux I__3694 (
            .O(N__17489),
            .I(N__17459));
    InMux I__3693 (
            .O(N__17488),
            .I(N__17459));
    InMux I__3692 (
            .O(N__17487),
            .I(N__17459));
    InMux I__3691 (
            .O(N__17486),
            .I(N__17459));
    InMux I__3690 (
            .O(N__17485),
            .I(N__17454));
    InMux I__3689 (
            .O(N__17484),
            .I(N__17454));
    Span4Mux_h I__3688 (
            .O(N__17477),
            .I(N__17451));
    InMux I__3687 (
            .O(N__17476),
            .I(N__17448));
    LocalMux I__3686 (
            .O(N__17473),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__3685 (
            .O(N__17468),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__3684 (
            .O(N__17459),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__3683 (
            .O(N__17454),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__3682 (
            .O(N__17451),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__3681 (
            .O(N__17448),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    InMux I__3680 (
            .O(N__17435),
            .I(N__17432));
    LocalMux I__3679 (
            .O(N__17432),
            .I(N__17429));
    Odrv4 I__3678 (
            .O(N__17429),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_41 ));
    InMux I__3677 (
            .O(N__17426),
            .I(N__17411));
    InMux I__3676 (
            .O(N__17425),
            .I(N__17411));
    InMux I__3675 (
            .O(N__17424),
            .I(N__17411));
    InMux I__3674 (
            .O(N__17423),
            .I(N__17406));
    InMux I__3673 (
            .O(N__17422),
            .I(N__17406));
    InMux I__3672 (
            .O(N__17421),
            .I(N__17403));
    InMux I__3671 (
            .O(N__17420),
            .I(N__17400));
    InMux I__3670 (
            .O(N__17419),
            .I(N__17397));
    CascadeMux I__3669 (
            .O(N__17418),
            .I(N__17392));
    LocalMux I__3668 (
            .O(N__17411),
            .I(N__17382));
    LocalMux I__3667 (
            .O(N__17406),
            .I(N__17382));
    LocalMux I__3666 (
            .O(N__17403),
            .I(N__17379));
    LocalMux I__3665 (
            .O(N__17400),
            .I(N__17374));
    LocalMux I__3664 (
            .O(N__17397),
            .I(N__17374));
    InMux I__3663 (
            .O(N__17396),
            .I(N__17369));
    InMux I__3662 (
            .O(N__17395),
            .I(N__17369));
    InMux I__3661 (
            .O(N__17392),
            .I(N__17366));
    InMux I__3660 (
            .O(N__17391),
            .I(N__17359));
    InMux I__3659 (
            .O(N__17390),
            .I(N__17359));
    InMux I__3658 (
            .O(N__17389),
            .I(N__17359));
    InMux I__3657 (
            .O(N__17388),
            .I(N__17354));
    InMux I__3656 (
            .O(N__17387),
            .I(N__17354));
    Span4Mux_h I__3655 (
            .O(N__17382),
            .I(N__17351));
    Span4Mux_v I__3654 (
            .O(N__17379),
            .I(N__17344));
    Span4Mux_v I__3653 (
            .O(N__17374),
            .I(N__17344));
    LocalMux I__3652 (
            .O(N__17369),
            .I(N__17344));
    LocalMux I__3651 (
            .O(N__17366),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__3650 (
            .O(N__17359),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__3649 (
            .O(N__17354),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__3648 (
            .O(N__17351),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__3647 (
            .O(N__17344),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    InMux I__3646 (
            .O(N__17333),
            .I(N__17329));
    InMux I__3645 (
            .O(N__17332),
            .I(N__17326));
    LocalMux I__3644 (
            .O(N__17329),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__3643 (
            .O(N__17326),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    CascadeMux I__3642 (
            .O(N__17321),
            .I(N__17317));
    InMux I__3641 (
            .O(N__17320),
            .I(N__17307));
    InMux I__3640 (
            .O(N__17317),
            .I(N__17307));
    InMux I__3639 (
            .O(N__17316),
            .I(N__17307));
    CascadeMux I__3638 (
            .O(N__17315),
            .I(N__17304));
    CascadeMux I__3637 (
            .O(N__17314),
            .I(N__17299));
    LocalMux I__3636 (
            .O(N__17307),
            .I(N__17293));
    InMux I__3635 (
            .O(N__17304),
            .I(N__17282));
    InMux I__3634 (
            .O(N__17303),
            .I(N__17282));
    InMux I__3633 (
            .O(N__17302),
            .I(N__17282));
    InMux I__3632 (
            .O(N__17299),
            .I(N__17282));
    InMux I__3631 (
            .O(N__17298),
            .I(N__17282));
    InMux I__3630 (
            .O(N__17297),
            .I(N__17276));
    InMux I__3629 (
            .O(N__17296),
            .I(N__17276));
    Span4Mux_h I__3628 (
            .O(N__17293),
            .I(N__17271));
    LocalMux I__3627 (
            .O(N__17282),
            .I(N__17271));
    InMux I__3626 (
            .O(N__17281),
            .I(N__17268));
    LocalMux I__3625 (
            .O(N__17276),
            .I(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5 ));
    Odrv4 I__3624 (
            .O(N__17271),
            .I(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5 ));
    LocalMux I__3623 (
            .O(N__17268),
            .I(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5 ));
    InMux I__3622 (
            .O(N__17261),
            .I(N__17258));
    LocalMux I__3621 (
            .O(N__17258),
            .I(N__17250));
    InMux I__3620 (
            .O(N__17257),
            .I(N__17243));
    InMux I__3619 (
            .O(N__17256),
            .I(N__17243));
    InMux I__3618 (
            .O(N__17255),
            .I(N__17240));
    InMux I__3617 (
            .O(N__17254),
            .I(N__17237));
    InMux I__3616 (
            .O(N__17253),
            .I(N__17234));
    Span4Mux_h I__3615 (
            .O(N__17250),
            .I(N__17231));
    InMux I__3614 (
            .O(N__17249),
            .I(N__17228));
    InMux I__3613 (
            .O(N__17248),
            .I(N__17225));
    LocalMux I__3612 (
            .O(N__17243),
            .I(N__17222));
    LocalMux I__3611 (
            .O(N__17240),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3610 (
            .O(N__17237),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3609 (
            .O(N__17234),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__3608 (
            .O(N__17231),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3607 (
            .O(N__17228),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__3606 (
            .O(N__17225),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__3605 (
            .O(N__17222),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    CascadeMux I__3604 (
            .O(N__17207),
            .I(N__17199));
    CascadeMux I__3603 (
            .O(N__17206),
            .I(N__17196));
    InMux I__3602 (
            .O(N__17205),
            .I(N__17189));
    InMux I__3601 (
            .O(N__17204),
            .I(N__17189));
    InMux I__3600 (
            .O(N__17203),
            .I(N__17189));
    InMux I__3599 (
            .O(N__17202),
            .I(N__17186));
    InMux I__3598 (
            .O(N__17199),
            .I(N__17181));
    InMux I__3597 (
            .O(N__17196),
            .I(N__17181));
    LocalMux I__3596 (
            .O(N__17189),
            .I(N__17175));
    LocalMux I__3595 (
            .O(N__17186),
            .I(N__17166));
    LocalMux I__3594 (
            .O(N__17181),
            .I(N__17166));
    InMux I__3593 (
            .O(N__17180),
            .I(N__17161));
    InMux I__3592 (
            .O(N__17179),
            .I(N__17161));
    InMux I__3591 (
            .O(N__17178),
            .I(N__17158));
    Span4Mux_h I__3590 (
            .O(N__17175),
            .I(N__17155));
    InMux I__3589 (
            .O(N__17174),
            .I(N__17152));
    InMux I__3588 (
            .O(N__17173),
            .I(N__17147));
    InMux I__3587 (
            .O(N__17172),
            .I(N__17147));
    InMux I__3586 (
            .O(N__17171),
            .I(N__17144));
    Span4Mux_h I__3585 (
            .O(N__17166),
            .I(N__17139));
    LocalMux I__3584 (
            .O(N__17161),
            .I(N__17139));
    LocalMux I__3583 (
            .O(N__17158),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__3582 (
            .O(N__17155),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__3581 (
            .O(N__17152),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__3580 (
            .O(N__17147),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__3579 (
            .O(N__17144),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__3578 (
            .O(N__17139),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__3577 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__3576 (
            .O(N__17123),
            .I(\uu2.mem0.G_11_0_0_a2_3_4 ));
    CascadeMux I__3575 (
            .O(N__17120),
            .I(N__17114));
    InMux I__3574 (
            .O(N__17119),
            .I(N__17111));
    InMux I__3573 (
            .O(N__17118),
            .I(N__17104));
    InMux I__3572 (
            .O(N__17117),
            .I(N__17104));
    InMux I__3571 (
            .O(N__17114),
            .I(N__17104));
    LocalMux I__3570 (
            .O(N__17111),
            .I(N__17099));
    LocalMux I__3569 (
            .O(N__17104),
            .I(N__17099));
    Span4Mux_s3_v I__3568 (
            .O(N__17099),
            .I(N__17096));
    Odrv4 I__3567 (
            .O(N__17096),
            .I(N_272_mux));
    CascadeMux I__3566 (
            .O(N__17093),
            .I(\uu2.mem0.G_11_0_0_a2_3_5_cascade_ ));
    InMux I__3565 (
            .O(N__17090),
            .I(N__17087));
    LocalMux I__3564 (
            .O(N__17087),
            .I(N__17083));
    InMux I__3563 (
            .O(N__17086),
            .I(N__17080));
    Span4Mux_s3_h I__3562 (
            .O(N__17083),
            .I(N__17077));
    LocalMux I__3561 (
            .O(N__17080),
            .I(N__17074));
    Span4Mux_h I__3560 (
            .O(N__17077),
            .I(N__17070));
    Span4Mux_h I__3559 (
            .O(N__17074),
            .I(N__17067));
    InMux I__3558 (
            .O(N__17073),
            .I(N__17064));
    Odrv4 I__3557 (
            .O(N__17070),
            .I(L3_tx_data_1));
    Odrv4 I__3556 (
            .O(N__17067),
            .I(L3_tx_data_1));
    LocalMux I__3555 (
            .O(N__17064),
            .I(L3_tx_data_1));
    InMux I__3554 (
            .O(N__17057),
            .I(N__17054));
    LocalMux I__3553 (
            .O(N__17054),
            .I(\uu2.mem0.G_11_0_0_0 ));
    InMux I__3552 (
            .O(N__17051),
            .I(N__17048));
    LocalMux I__3551 (
            .O(N__17048),
            .I(N__17045));
    Span4Mux_h I__3550 (
            .O(N__17045),
            .I(N__17042));
    Odrv4 I__3549 (
            .O(N__17042),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_1 ));
    InMux I__3548 (
            .O(N__17039),
            .I(N__17036));
    LocalMux I__3547 (
            .O(N__17036),
            .I(N__17033));
    Span4Mux_v I__3546 (
            .O(N__17033),
            .I(N__17030));
    Odrv4 I__3545 (
            .O(N__17030),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_5 ));
    InMux I__3544 (
            .O(N__17027),
            .I(N__17024));
    LocalMux I__3543 (
            .O(N__17024),
            .I(N__17021));
    Span4Mux_h I__3542 (
            .O(N__17021),
            .I(N__17018));
    Odrv4 I__3541 (
            .O(N__17018),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_4 ));
    InMux I__3540 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__3539 (
            .O(N__17012),
            .I(N__17009));
    Span4Mux_h I__3538 (
            .O(N__17009),
            .I(N__17006));
    Odrv4 I__3537 (
            .O(N__17006),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_2 ));
    InMux I__3536 (
            .O(N__17003),
            .I(N__17000));
    LocalMux I__3535 (
            .O(N__17000),
            .I(\uu2.bitmapZ0Z_212 ));
    CascadeMux I__3534 (
            .O(N__16997),
            .I(N__16994));
    InMux I__3533 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__3532 (
            .O(N__16991),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__3531 (
            .O(N__16988),
            .I(N__16985));
    LocalMux I__3530 (
            .O(N__16985),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__3529 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__3528 (
            .O(N__16979),
            .I(\uu2.bitmapZ0Z_84 ));
    CascadeMux I__3527 (
            .O(N__16976),
            .I(\uu2.bitmap_pmux_17_ns_1_cascade_ ));
    CascadeMux I__3526 (
            .O(N__16973),
            .I(N__16963));
    CascadeMux I__3525 (
            .O(N__16972),
            .I(N__16958));
    CascadeMux I__3524 (
            .O(N__16971),
            .I(N__16954));
    InMux I__3523 (
            .O(N__16970),
            .I(N__16951));
    InMux I__3522 (
            .O(N__16969),
            .I(N__16946));
    InMux I__3521 (
            .O(N__16968),
            .I(N__16943));
    InMux I__3520 (
            .O(N__16967),
            .I(N__16940));
    CascadeMux I__3519 (
            .O(N__16966),
            .I(N__16937));
    InMux I__3518 (
            .O(N__16963),
            .I(N__16932));
    InMux I__3517 (
            .O(N__16962),
            .I(N__16932));
    InMux I__3516 (
            .O(N__16961),
            .I(N__16923));
    InMux I__3515 (
            .O(N__16958),
            .I(N__16923));
    InMux I__3514 (
            .O(N__16957),
            .I(N__16923));
    InMux I__3513 (
            .O(N__16954),
            .I(N__16923));
    LocalMux I__3512 (
            .O(N__16951),
            .I(N__16920));
    InMux I__3511 (
            .O(N__16950),
            .I(N__16917));
    InMux I__3510 (
            .O(N__16949),
            .I(N__16914));
    LocalMux I__3509 (
            .O(N__16946),
            .I(N__16909));
    LocalMux I__3508 (
            .O(N__16943),
            .I(N__16909));
    LocalMux I__3507 (
            .O(N__16940),
            .I(N__16906));
    InMux I__3506 (
            .O(N__16937),
            .I(N__16903));
    LocalMux I__3505 (
            .O(N__16932),
            .I(N__16900));
    LocalMux I__3504 (
            .O(N__16923),
            .I(N__16891));
    Span4Mux_h I__3503 (
            .O(N__16920),
            .I(N__16891));
    LocalMux I__3502 (
            .O(N__16917),
            .I(N__16891));
    LocalMux I__3501 (
            .O(N__16914),
            .I(N__16891));
    Span4Mux_v I__3500 (
            .O(N__16909),
            .I(N__16886));
    Span4Mux_v I__3499 (
            .O(N__16906),
            .I(N__16886));
    LocalMux I__3498 (
            .O(N__16903),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv12 I__3497 (
            .O(N__16900),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3496 (
            .O(N__16891),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3495 (
            .O(N__16886),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    CascadeMux I__3494 (
            .O(N__16877),
            .I(\Lab_UT.dictrl.g0_8Z0Z_3_cascade_ ));
    CascadeMux I__3493 (
            .O(N__16874),
            .I(N__16871));
    InMux I__3492 (
            .O(N__16871),
            .I(N__16868));
    LocalMux I__3491 (
            .O(N__16868),
            .I(N__16865));
    Odrv4 I__3490 (
            .O(N__16865),
            .I(\Lab_UT.dictrl.g2_1_3 ));
    InMux I__3489 (
            .O(N__16862),
            .I(N__16854));
    InMux I__3488 (
            .O(N__16861),
            .I(N__16854));
    InMux I__3487 (
            .O(N__16860),
            .I(N__16851));
    InMux I__3486 (
            .O(N__16859),
            .I(N__16848));
    LocalMux I__3485 (
            .O(N__16854),
            .I(N__16843));
    LocalMux I__3484 (
            .O(N__16851),
            .I(N__16843));
    LocalMux I__3483 (
            .O(N__16848),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__3482 (
            .O(N__16843),
            .I(bu_rx_data_1_rep1));
    InMux I__3481 (
            .O(N__16838),
            .I(N__16835));
    LocalMux I__3480 (
            .O(N__16835),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_28 ));
    InMux I__3479 (
            .O(N__16832),
            .I(N__16829));
    LocalMux I__3478 (
            .O(N__16829),
            .I(\uu2.mem0.N_44 ));
    CascadeMux I__3477 (
            .O(N__16826),
            .I(\uu2.mem0.N_41_cascade_ ));
    InMux I__3476 (
            .O(N__16823),
            .I(N__16820));
    LocalMux I__3475 (
            .O(N__16820),
            .I(N__16817));
    Span4Mux_h I__3474 (
            .O(N__16817),
            .I(N__16814));
    Odrv4 I__3473 (
            .O(N__16814),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__3472 (
            .O(N__16811),
            .I(N__16805));
    InMux I__3471 (
            .O(N__16810),
            .I(N__16805));
    LocalMux I__3470 (
            .O(N__16805),
            .I(N__16802));
    Span4Mux_h I__3469 (
            .O(N__16802),
            .I(N__16798));
    InMux I__3468 (
            .O(N__16801),
            .I(N__16795));
    Odrv4 I__3467 (
            .O(N__16798),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    LocalMux I__3466 (
            .O(N__16795),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    CascadeMux I__3465 (
            .O(N__16790),
            .I(\uu2.mem0.N_24_i_cascade_ ));
    InMux I__3464 (
            .O(N__16787),
            .I(N__16782));
    InMux I__3463 (
            .O(N__16786),
            .I(N__16779));
    InMux I__3462 (
            .O(N__16785),
            .I(N__16776));
    LocalMux I__3461 (
            .O(N__16782),
            .I(N__16773));
    LocalMux I__3460 (
            .O(N__16779),
            .I(\uu2.N_406 ));
    LocalMux I__3459 (
            .O(N__16776),
            .I(\uu2.N_406 ));
    Odrv12 I__3458 (
            .O(N__16773),
            .I(\uu2.N_406 ));
    InMux I__3457 (
            .O(N__16766),
            .I(N__16763));
    LocalMux I__3456 (
            .O(N__16763),
            .I(\uu2.mem0.N_45 ));
    InMux I__3455 (
            .O(N__16760),
            .I(N__16757));
    LocalMux I__3454 (
            .O(N__16757),
            .I(N__16754));
    Odrv12 I__3453 (
            .O(N__16754),
            .I(\Lab_UT.dictrl.next_alarmstate4Z0Z_3 ));
    InMux I__3452 (
            .O(N__16751),
            .I(N__16748));
    LocalMux I__3451 (
            .O(N__16748),
            .I(N__16745));
    Odrv4 I__3450 (
            .O(N__16745),
            .I(\Lab_UT.dictrl.next_alarmstate4Z0Z_0 ));
    InMux I__3449 (
            .O(N__16742),
            .I(N__16739));
    LocalMux I__3448 (
            .O(N__16739),
            .I(\Lab_UT.dictrl.g2_1_2 ));
    CascadeMux I__3447 (
            .O(N__16736),
            .I(\Lab_UT.dictrl.g1_5_1_cascade_ ));
    InMux I__3446 (
            .O(N__16733),
            .I(N__16730));
    LocalMux I__3445 (
            .O(N__16730),
            .I(\Lab_UT.dictrl.g2_3 ));
    InMux I__3444 (
            .O(N__16727),
            .I(N__16724));
    LocalMux I__3443 (
            .O(N__16724),
            .I(\Lab_UT.dictrl.g0Z0Z_1 ));
    CascadeMux I__3442 (
            .O(N__16721),
            .I(\Lab_UT.dictrl.g0_3_cascade_ ));
    InMux I__3441 (
            .O(N__16718),
            .I(N__16708));
    InMux I__3440 (
            .O(N__16717),
            .I(N__16703));
    InMux I__3439 (
            .O(N__16716),
            .I(N__16703));
    InMux I__3438 (
            .O(N__16715),
            .I(N__16696));
    InMux I__3437 (
            .O(N__16714),
            .I(N__16696));
    InMux I__3436 (
            .O(N__16713),
            .I(N__16696));
    InMux I__3435 (
            .O(N__16712),
            .I(N__16691));
    InMux I__3434 (
            .O(N__16711),
            .I(N__16691));
    LocalMux I__3433 (
            .O(N__16708),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3432 (
            .O(N__16703),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3431 (
            .O(N__16696),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3430 (
            .O(N__16691),
            .I(bu_rx_data_5_rep1));
    InMux I__3429 (
            .O(N__16682),
            .I(N__16676));
    InMux I__3428 (
            .O(N__16681),
            .I(N__16676));
    LocalMux I__3427 (
            .O(N__16676),
            .I(N__16673));
    Odrv4 I__3426 (
            .O(N__16673),
            .I(\Lab_UT.dictrl.next_state12_0 ));
    CascadeMux I__3425 (
            .O(N__16670),
            .I(N__16665));
    InMux I__3424 (
            .O(N__16669),
            .I(N__16660));
    CascadeMux I__3423 (
            .O(N__16668),
            .I(N__16656));
    InMux I__3422 (
            .O(N__16665),
            .I(N__16647));
    InMux I__3421 (
            .O(N__16664),
            .I(N__16647));
    InMux I__3420 (
            .O(N__16663),
            .I(N__16647));
    LocalMux I__3419 (
            .O(N__16660),
            .I(N__16644));
    InMux I__3418 (
            .O(N__16659),
            .I(N__16637));
    InMux I__3417 (
            .O(N__16656),
            .I(N__16637));
    InMux I__3416 (
            .O(N__16655),
            .I(N__16637));
    InMux I__3415 (
            .O(N__16654),
            .I(N__16634));
    LocalMux I__3414 (
            .O(N__16647),
            .I(N__16631));
    Odrv4 I__3413 (
            .O(N__16644),
            .I(bu_rx_data_6_rep1));
    LocalMux I__3412 (
            .O(N__16637),
            .I(bu_rx_data_6_rep1));
    LocalMux I__3411 (
            .O(N__16634),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__3410 (
            .O(N__16631),
            .I(bu_rx_data_6_rep1));
    CascadeMux I__3409 (
            .O(N__16622),
            .I(N__16619));
    InMux I__3408 (
            .O(N__16619),
            .I(N__16616));
    LocalMux I__3407 (
            .O(N__16616),
            .I(\Lab_UT.dictrl.g0_0_0_o4_0 ));
    CascadeMux I__3406 (
            .O(N__16613),
            .I(\Lab_UT.dictrl.N_3_0_cascade_ ));
    InMux I__3405 (
            .O(N__16610),
            .I(N__16607));
    LocalMux I__3404 (
            .O(N__16607),
            .I(\Lab_UT.dictrl.g0_0_0_a3_2_0 ));
    InMux I__3403 (
            .O(N__16604),
            .I(N__16601));
    LocalMux I__3402 (
            .O(N__16601),
            .I(N__16598));
    Odrv4 I__3401 (
            .O(N__16598),
            .I(\Lab_UT.dictrl.g0_0_i_o4_0 ));
    InMux I__3400 (
            .O(N__16595),
            .I(N__16584));
    InMux I__3399 (
            .O(N__16594),
            .I(N__16584));
    InMux I__3398 (
            .O(N__16593),
            .I(N__16584));
    InMux I__3397 (
            .O(N__16592),
            .I(N__16579));
    InMux I__3396 (
            .O(N__16591),
            .I(N__16579));
    LocalMux I__3395 (
            .O(N__16584),
            .I(N__16573));
    LocalMux I__3394 (
            .O(N__16579),
            .I(N__16570));
    InMux I__3393 (
            .O(N__16578),
            .I(N__16563));
    InMux I__3392 (
            .O(N__16577),
            .I(N__16563));
    InMux I__3391 (
            .O(N__16576),
            .I(N__16563));
    Odrv4 I__3390 (
            .O(N__16573),
            .I(\Lab_UT.dictrl.g0_1Z0Z_2 ));
    Odrv4 I__3389 (
            .O(N__16570),
            .I(\Lab_UT.dictrl.g0_1Z0Z_2 ));
    LocalMux I__3388 (
            .O(N__16563),
            .I(\Lab_UT.dictrl.g0_1Z0Z_2 ));
    InMux I__3387 (
            .O(N__16556),
            .I(N__16553));
    LocalMux I__3386 (
            .O(N__16553),
            .I(\Lab_UT.dictrl.next_state18_0 ));
    CascadeMux I__3385 (
            .O(N__16550),
            .I(\Lab_UT.dictrl.next_state18_0_cascade_ ));
    CascadeMux I__3384 (
            .O(N__16547),
            .I(\Lab_UT.dictrl.g2_0_0_cascade_ ));
    InMux I__3383 (
            .O(N__16544),
            .I(N__16541));
    LocalMux I__3382 (
            .O(N__16541),
            .I(\Lab_UT.dictrl.N_7_0 ));
    InMux I__3381 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__3380 (
            .O(N__16535),
            .I(N__16532));
    Odrv12 I__3379 (
            .O(N__16532),
            .I(\Lab_UT.dictrl.N_11 ));
    InMux I__3378 (
            .O(N__16529),
            .I(N__16526));
    LocalMux I__3377 (
            .O(N__16526),
            .I(\Lab_UT.dictrl.g2_2_0 ));
    InMux I__3376 (
            .O(N__16523),
            .I(N__16520));
    LocalMux I__3375 (
            .O(N__16520),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_3_0 ));
    InMux I__3374 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__3373 (
            .O(N__16514),
            .I(N__16511));
    Odrv4 I__3372 (
            .O(N__16511),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_4 ));
    InMux I__3371 (
            .O(N__16508),
            .I(N__16505));
    LocalMux I__3370 (
            .O(N__16505),
            .I(N__16502));
    Sp12to4 I__3369 (
            .O(N__16502),
            .I(N__16499));
    Odrv12 I__3368 (
            .O(N__16499),
            .I(\Lab_UT.dictrl.N_9_0 ));
    CascadeMux I__3367 (
            .O(N__16496),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_ ));
    InMux I__3366 (
            .O(N__16493),
            .I(N__16483));
    InMux I__3365 (
            .O(N__16492),
            .I(N__16483));
    InMux I__3364 (
            .O(N__16491),
            .I(N__16479));
    InMux I__3363 (
            .O(N__16490),
            .I(N__16476));
    InMux I__3362 (
            .O(N__16489),
            .I(N__16471));
    InMux I__3361 (
            .O(N__16488),
            .I(N__16468));
    LocalMux I__3360 (
            .O(N__16483),
            .I(N__16465));
    InMux I__3359 (
            .O(N__16482),
            .I(N__16462));
    LocalMux I__3358 (
            .O(N__16479),
            .I(N__16459));
    LocalMux I__3357 (
            .O(N__16476),
            .I(N__16456));
    InMux I__3356 (
            .O(N__16475),
            .I(N__16451));
    InMux I__3355 (
            .O(N__16474),
            .I(N__16451));
    LocalMux I__3354 (
            .O(N__16471),
            .I(N__16447));
    LocalMux I__3353 (
            .O(N__16468),
            .I(N__16440));
    Span4Mux_v I__3352 (
            .O(N__16465),
            .I(N__16440));
    LocalMux I__3351 (
            .O(N__16462),
            .I(N__16440));
    Span4Mux_h I__3350 (
            .O(N__16459),
            .I(N__16435));
    Span4Mux_v I__3349 (
            .O(N__16456),
            .I(N__16435));
    LocalMux I__3348 (
            .O(N__16451),
            .I(N__16432));
    InMux I__3347 (
            .O(N__16450),
            .I(N__16429));
    Span4Mux_h I__3346 (
            .O(N__16447),
            .I(N__16424));
    Span4Mux_h I__3345 (
            .O(N__16440),
            .I(N__16424));
    Odrv4 I__3344 (
            .O(N__16435),
            .I(bu_rx_data_0));
    Odrv12 I__3343 (
            .O(N__16432),
            .I(bu_rx_data_0));
    LocalMux I__3342 (
            .O(N__16429),
            .I(bu_rx_data_0));
    Odrv4 I__3341 (
            .O(N__16424),
            .I(bu_rx_data_0));
    InMux I__3340 (
            .O(N__16415),
            .I(N__16409));
    InMux I__3339 (
            .O(N__16414),
            .I(N__16409));
    LocalMux I__3338 (
            .O(N__16409),
            .I(N__16406));
    Span4Mux_h I__3337 (
            .O(N__16406),
            .I(N__16403));
    Odrv4 I__3336 (
            .O(N__16403),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z4 ));
    CascadeMux I__3335 (
            .O(N__16400),
            .I(\Lab_UT.dictrl.N_5_cascade_ ));
    InMux I__3334 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__3333 (
            .O(N__16394),
            .I(\Lab_UT.dictrl.N_10_0 ));
    CascadeMux I__3332 (
            .O(N__16391),
            .I(N__16386));
    CascadeMux I__3331 (
            .O(N__16390),
            .I(N__16382));
    InMux I__3330 (
            .O(N__16389),
            .I(N__16375));
    InMux I__3329 (
            .O(N__16386),
            .I(N__16375));
    InMux I__3328 (
            .O(N__16385),
            .I(N__16375));
    InMux I__3327 (
            .O(N__16382),
            .I(N__16372));
    LocalMux I__3326 (
            .O(N__16375),
            .I(N__16369));
    LocalMux I__3325 (
            .O(N__16372),
            .I(N__16366));
    Span12Mux_s7_h I__3324 (
            .O(N__16369),
            .I(N__16363));
    Span4Mux_v I__3323 (
            .O(N__16366),
            .I(N__16360));
    Odrv12 I__3322 (
            .O(N__16363),
            .I(\Lab_UT.dicRun_2 ));
    Odrv4 I__3321 (
            .O(N__16360),
            .I(\Lab_UT.dicRun_2 ));
    InMux I__3320 (
            .O(N__16355),
            .I(N__16352));
    LocalMux I__3319 (
            .O(N__16352),
            .I(\Lab_UT.didp.ce_9_0_0 ));
    CascadeMux I__3318 (
            .O(N__16349),
            .I(\Lab_UT.dicRun_2_cascade_ ));
    InMux I__3317 (
            .O(N__16346),
            .I(N__16341));
    InMux I__3316 (
            .O(N__16345),
            .I(N__16338));
    InMux I__3315 (
            .O(N__16344),
            .I(N__16331));
    LocalMux I__3314 (
            .O(N__16341),
            .I(N__16326));
    LocalMux I__3313 (
            .O(N__16338),
            .I(N__16326));
    InMux I__3312 (
            .O(N__16337),
            .I(N__16323));
    InMux I__3311 (
            .O(N__16336),
            .I(N__16318));
    InMux I__3310 (
            .O(N__16335),
            .I(N__16318));
    InMux I__3309 (
            .O(N__16334),
            .I(N__16313));
    LocalMux I__3308 (
            .O(N__16331),
            .I(N__16310));
    Span4Mux_v I__3307 (
            .O(N__16326),
            .I(N__16305));
    LocalMux I__3306 (
            .O(N__16323),
            .I(N__16305));
    LocalMux I__3305 (
            .O(N__16318),
            .I(N__16302));
    InMux I__3304 (
            .O(N__16317),
            .I(N__16294));
    InMux I__3303 (
            .O(N__16316),
            .I(N__16294));
    LocalMux I__3302 (
            .O(N__16313),
            .I(N__16289));
    Span4Mux_v I__3301 (
            .O(N__16310),
            .I(N__16286));
    Span4Mux_h I__3300 (
            .O(N__16305),
            .I(N__16281));
    Span4Mux_h I__3299 (
            .O(N__16302),
            .I(N__16281));
    InMux I__3298 (
            .O(N__16301),
            .I(N__16274));
    InMux I__3297 (
            .O(N__16300),
            .I(N__16274));
    InMux I__3296 (
            .O(N__16299),
            .I(N__16274));
    LocalMux I__3295 (
            .O(N__16294),
            .I(N__16271));
    InMux I__3294 (
            .O(N__16293),
            .I(N__16266));
    InMux I__3293 (
            .O(N__16292),
            .I(N__16266));
    Span4Mux_v I__3292 (
            .O(N__16289),
            .I(N__16259));
    Span4Mux_h I__3291 (
            .O(N__16286),
            .I(N__16259));
    Span4Mux_v I__3290 (
            .O(N__16281),
            .I(N__16259));
    LocalMux I__3289 (
            .O(N__16274),
            .I(oneSecStrb));
    Odrv4 I__3288 (
            .O(N__16271),
            .I(oneSecStrb));
    LocalMux I__3287 (
            .O(N__16266),
            .I(oneSecStrb));
    Odrv4 I__3286 (
            .O(N__16259),
            .I(oneSecStrb));
    InMux I__3285 (
            .O(N__16250),
            .I(N__16240));
    InMux I__3284 (
            .O(N__16249),
            .I(N__16240));
    InMux I__3283 (
            .O(N__16248),
            .I(N__16240));
    InMux I__3282 (
            .O(N__16247),
            .I(N__16237));
    LocalMux I__3281 (
            .O(N__16240),
            .I(N__16234));
    LocalMux I__3280 (
            .O(N__16237),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    Odrv4 I__3279 (
            .O(N__16234),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__3278 (
            .O(N__16229),
            .I(N__16226));
    LocalMux I__3277 (
            .O(N__16226),
            .I(\Lab_UT.dictrl.N_11_0 ));
    CascadeMux I__3276 (
            .O(N__16223),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_ ));
    InMux I__3275 (
            .O(N__16220),
            .I(N__16217));
    LocalMux I__3274 (
            .O(N__16217),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_1 ));
    InMux I__3273 (
            .O(N__16214),
            .I(N__16211));
    LocalMux I__3272 (
            .O(N__16211),
            .I(\Lab_UT.dictrl.g0_0_i_a3_3_1 ));
    InMux I__3271 (
            .O(N__16208),
            .I(N__16205));
    LocalMux I__3270 (
            .O(N__16205),
            .I(\Lab_UT.bcd2segment3.segment_0Z0Z_2 ));
    InMux I__3269 (
            .O(N__16202),
            .I(N__16199));
    LocalMux I__3268 (
            .O(N__16199),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_4 ));
    InMux I__3267 (
            .O(N__16196),
            .I(N__16193));
    LocalMux I__3266 (
            .O(N__16193),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_6 ));
    InMux I__3265 (
            .O(N__16190),
            .I(N__16187));
    LocalMux I__3264 (
            .O(N__16187),
            .I(N__16184));
    Odrv12 I__3263 (
            .O(N__16184),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__3262 (
            .O(N__16181),
            .I(N__16178));
    LocalMux I__3261 (
            .O(N__16178),
            .I(\Lab_UT.bcd2segment3.segment_0Z0Z_1 ));
    InMux I__3260 (
            .O(N__16175),
            .I(N__16172));
    LocalMux I__3259 (
            .O(N__16172),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_5 ));
    InMux I__3258 (
            .O(N__16169),
            .I(N__16166));
    LocalMux I__3257 (
            .O(N__16166),
            .I(N__16163));
    Odrv4 I__3256 (
            .O(N__16163),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__3255 (
            .O(N__16160),
            .I(N__16157));
    LocalMux I__3254 (
            .O(N__16157),
            .I(N__16154));
    Span4Mux_h I__3253 (
            .O(N__16154),
            .I(N__16151));
    Odrv4 I__3252 (
            .O(N__16151),
            .I(\Lab_UT.LdASones ));
    CascadeMux I__3251 (
            .O(N__16148),
            .I(\Lab_UT.LdASones_cascade_ ));
    InMux I__3250 (
            .O(N__16145),
            .I(N__16142));
    LocalMux I__3249 (
            .O(N__16142),
            .I(N__16139));
    Span4Mux_v I__3248 (
            .O(N__16139),
            .I(N__16136));
    Odrv4 I__3247 (
            .O(N__16136),
            .I(\Lab_UT.LdSones_i_3 ));
    InMux I__3246 (
            .O(N__16133),
            .I(N__16130));
    LocalMux I__3245 (
            .O(N__16130),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__3244 (
            .O(N__16127),
            .I(N__16122));
    CascadeMux I__3243 (
            .O(N__16126),
            .I(N__16110));
    InMux I__3242 (
            .O(N__16125),
            .I(N__16106));
    LocalMux I__3241 (
            .O(N__16122),
            .I(N__16103));
    InMux I__3240 (
            .O(N__16121),
            .I(N__16100));
    InMux I__3239 (
            .O(N__16120),
            .I(N__16095));
    InMux I__3238 (
            .O(N__16119),
            .I(N__16095));
    InMux I__3237 (
            .O(N__16118),
            .I(N__16090));
    InMux I__3236 (
            .O(N__16117),
            .I(N__16090));
    InMux I__3235 (
            .O(N__16116),
            .I(N__16083));
    InMux I__3234 (
            .O(N__16115),
            .I(N__16083));
    InMux I__3233 (
            .O(N__16114),
            .I(N__16083));
    InMux I__3232 (
            .O(N__16113),
            .I(N__16076));
    InMux I__3231 (
            .O(N__16110),
            .I(N__16076));
    InMux I__3230 (
            .O(N__16109),
            .I(N__16076));
    LocalMux I__3229 (
            .O(N__16106),
            .I(N__16073));
    Odrv4 I__3228 (
            .O(N__16103),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3227 (
            .O(N__16100),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3226 (
            .O(N__16095),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3225 (
            .O(N__16090),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3224 (
            .O(N__16083),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__3223 (
            .O(N__16076),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__3222 (
            .O(N__16073),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CascadeMux I__3221 (
            .O(N__16058),
            .I(\uu2.N_98_cascade_ ));
    InMux I__3220 (
            .O(N__16055),
            .I(N__16049));
    InMux I__3219 (
            .O(N__16054),
            .I(N__16049));
    LocalMux I__3218 (
            .O(N__16049),
            .I(\uu2.bitmap_RNI04AD1Z0Z_314 ));
    CascadeMux I__3217 (
            .O(N__16046),
            .I(N__16043));
    InMux I__3216 (
            .O(N__16043),
            .I(N__16036));
    InMux I__3215 (
            .O(N__16042),
            .I(N__16033));
    InMux I__3214 (
            .O(N__16041),
            .I(N__16028));
    InMux I__3213 (
            .O(N__16040),
            .I(N__16028));
    InMux I__3212 (
            .O(N__16039),
            .I(N__16025));
    LocalMux I__3211 (
            .O(N__16036),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__3210 (
            .O(N__16033),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__3209 (
            .O(N__16028),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__3208 (
            .O(N__16025),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__3207 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__3206 (
            .O(N__16013),
            .I(\uu2.bitmapZ0Z_180 ));
    InMux I__3205 (
            .O(N__16010),
            .I(N__16004));
    InMux I__3204 (
            .O(N__16009),
            .I(N__16004));
    LocalMux I__3203 (
            .O(N__16004),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__3202 (
            .O(N__16001),
            .I(N__15998));
    LocalMux I__3201 (
            .O(N__15998),
            .I(\uu2.N_383 ));
    CascadeMux I__3200 (
            .O(N__15995),
            .I(N__15989));
    InMux I__3199 (
            .O(N__15994),
            .I(N__15974));
    InMux I__3198 (
            .O(N__15993),
            .I(N__15969));
    InMux I__3197 (
            .O(N__15992),
            .I(N__15969));
    InMux I__3196 (
            .O(N__15989),
            .I(N__15962));
    InMux I__3195 (
            .O(N__15988),
            .I(N__15962));
    InMux I__3194 (
            .O(N__15987),
            .I(N__15962));
    InMux I__3193 (
            .O(N__15986),
            .I(N__15958));
    InMux I__3192 (
            .O(N__15985),
            .I(N__15955));
    InMux I__3191 (
            .O(N__15984),
            .I(N__15952));
    CascadeMux I__3190 (
            .O(N__15983),
            .I(N__15949));
    CascadeMux I__3189 (
            .O(N__15982),
            .I(N__15944));
    InMux I__3188 (
            .O(N__15981),
            .I(N__15933));
    InMux I__3187 (
            .O(N__15980),
            .I(N__15933));
    InMux I__3186 (
            .O(N__15979),
            .I(N__15933));
    InMux I__3185 (
            .O(N__15978),
            .I(N__15933));
    InMux I__3184 (
            .O(N__15977),
            .I(N__15933));
    LocalMux I__3183 (
            .O(N__15974),
            .I(N__15930));
    LocalMux I__3182 (
            .O(N__15969),
            .I(N__15926));
    LocalMux I__3181 (
            .O(N__15962),
            .I(N__15923));
    InMux I__3180 (
            .O(N__15961),
            .I(N__15920));
    LocalMux I__3179 (
            .O(N__15958),
            .I(N__15917));
    LocalMux I__3178 (
            .O(N__15955),
            .I(N__15912));
    LocalMux I__3177 (
            .O(N__15952),
            .I(N__15912));
    InMux I__3176 (
            .O(N__15949),
            .I(N__15903));
    InMux I__3175 (
            .O(N__15948),
            .I(N__15903));
    InMux I__3174 (
            .O(N__15947),
            .I(N__15903));
    InMux I__3173 (
            .O(N__15944),
            .I(N__15903));
    LocalMux I__3172 (
            .O(N__15933),
            .I(N__15898));
    Span4Mux_s2_v I__3171 (
            .O(N__15930),
            .I(N__15898));
    InMux I__3170 (
            .O(N__15929),
            .I(N__15895));
    Span4Mux_h I__3169 (
            .O(N__15926),
            .I(N__15892));
    Span4Mux_h I__3168 (
            .O(N__15923),
            .I(N__15889));
    LocalMux I__3167 (
            .O(N__15920),
            .I(N__15886));
    Span4Mux_h I__3166 (
            .O(N__15917),
            .I(N__15881));
    Span4Mux_h I__3165 (
            .O(N__15912),
            .I(N__15881));
    LocalMux I__3164 (
            .O(N__15903),
            .I(N__15876));
    Span4Mux_h I__3163 (
            .O(N__15898),
            .I(N__15876));
    LocalMux I__3162 (
            .O(N__15895),
            .I(N__15873));
    Odrv4 I__3161 (
            .O(N__15892),
            .I(L3_tx_data_rdy));
    Odrv4 I__3160 (
            .O(N__15889),
            .I(L3_tx_data_rdy));
    Odrv4 I__3159 (
            .O(N__15886),
            .I(L3_tx_data_rdy));
    Odrv4 I__3158 (
            .O(N__15881),
            .I(L3_tx_data_rdy));
    Odrv4 I__3157 (
            .O(N__15876),
            .I(L3_tx_data_rdy));
    Odrv12 I__3156 (
            .O(N__15873),
            .I(L3_tx_data_rdy));
    InMux I__3155 (
            .O(N__15860),
            .I(N__15845));
    InMux I__3154 (
            .O(N__15859),
            .I(N__15845));
    InMux I__3153 (
            .O(N__15858),
            .I(N__15845));
    InMux I__3152 (
            .O(N__15857),
            .I(N__15845));
    CascadeMux I__3151 (
            .O(N__15856),
            .I(N__15841));
    InMux I__3150 (
            .O(N__15855),
            .I(N__15832));
    InMux I__3149 (
            .O(N__15854),
            .I(N__15829));
    LocalMux I__3148 (
            .O(N__15845),
            .I(N__15822));
    InMux I__3147 (
            .O(N__15844),
            .I(N__15815));
    InMux I__3146 (
            .O(N__15841),
            .I(N__15815));
    InMux I__3145 (
            .O(N__15840),
            .I(N__15815));
    InMux I__3144 (
            .O(N__15839),
            .I(N__15804));
    InMux I__3143 (
            .O(N__15838),
            .I(N__15804));
    InMux I__3142 (
            .O(N__15837),
            .I(N__15804));
    InMux I__3141 (
            .O(N__15836),
            .I(N__15804));
    InMux I__3140 (
            .O(N__15835),
            .I(N__15804));
    LocalMux I__3139 (
            .O(N__15832),
            .I(N__15800));
    LocalMux I__3138 (
            .O(N__15829),
            .I(N__15797));
    InMux I__3137 (
            .O(N__15828),
            .I(N__15794));
    InMux I__3136 (
            .O(N__15827),
            .I(N__15789));
    InMux I__3135 (
            .O(N__15826),
            .I(N__15789));
    InMux I__3134 (
            .O(N__15825),
            .I(N__15786));
    Span4Mux_h I__3133 (
            .O(N__15822),
            .I(N__15783));
    LocalMux I__3132 (
            .O(N__15815),
            .I(N__15778));
    LocalMux I__3131 (
            .O(N__15804),
            .I(N__15778));
    InMux I__3130 (
            .O(N__15803),
            .I(N__15775));
    Span4Mux_h I__3129 (
            .O(N__15800),
            .I(N__15770));
    Span4Mux_s2_v I__3128 (
            .O(N__15797),
            .I(N__15770));
    LocalMux I__3127 (
            .O(N__15794),
            .I(uu2_un1_w_user_cr_0));
    LocalMux I__3126 (
            .O(N__15789),
            .I(uu2_un1_w_user_cr_0));
    LocalMux I__3125 (
            .O(N__15786),
            .I(uu2_un1_w_user_cr_0));
    Odrv4 I__3124 (
            .O(N__15783),
            .I(uu2_un1_w_user_cr_0));
    Odrv4 I__3123 (
            .O(N__15778),
            .I(uu2_un1_w_user_cr_0));
    LocalMux I__3122 (
            .O(N__15775),
            .I(uu2_un1_w_user_cr_0));
    Odrv4 I__3121 (
            .O(N__15770),
            .I(uu2_un1_w_user_cr_0));
    InMux I__3120 (
            .O(N__15755),
            .I(N__15749));
    InMux I__3119 (
            .O(N__15754),
            .I(N__15749));
    LocalMux I__3118 (
            .O(N__15749),
            .I(N__15745));
    CascadeMux I__3117 (
            .O(N__15748),
            .I(N__15742));
    Span4Mux_h I__3116 (
            .O(N__15745),
            .I(N__15738));
    InMux I__3115 (
            .O(N__15742),
            .I(N__15735));
    InMux I__3114 (
            .O(N__15741),
            .I(N__15732));
    Odrv4 I__3113 (
            .O(N__15738),
            .I(\uu2.N_57 ));
    LocalMux I__3112 (
            .O(N__15735),
            .I(\uu2.N_57 ));
    LocalMux I__3111 (
            .O(N__15732),
            .I(\uu2.N_57 ));
    CascadeMux I__3110 (
            .O(N__15725),
            .I(N__15719));
    InMux I__3109 (
            .O(N__15724),
            .I(N__15709));
    InMux I__3108 (
            .O(N__15723),
            .I(N__15709));
    InMux I__3107 (
            .O(N__15722),
            .I(N__15709));
    InMux I__3106 (
            .O(N__15719),
            .I(N__15709));
    CascadeMux I__3105 (
            .O(N__15718),
            .I(N__15706));
    LocalMux I__3104 (
            .O(N__15709),
            .I(N__15703));
    InMux I__3103 (
            .O(N__15706),
            .I(N__15700));
    Span4Mux_h I__3102 (
            .O(N__15703),
            .I(N__15697));
    LocalMux I__3101 (
            .O(N__15700),
            .I(\uu2.N_38 ));
    Odrv4 I__3100 (
            .O(N__15697),
            .I(\uu2.N_38 ));
    CascadeMux I__3099 (
            .O(N__15692),
            .I(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_ ));
    CascadeMux I__3098 (
            .O(N__15689),
            .I(N__15686));
    InMux I__3097 (
            .O(N__15686),
            .I(N__15682));
    CascadeMux I__3096 (
            .O(N__15685),
            .I(N__15675));
    LocalMux I__3095 (
            .O(N__15682),
            .I(N__15672));
    InMux I__3094 (
            .O(N__15681),
            .I(N__15668));
    InMux I__3093 (
            .O(N__15680),
            .I(N__15659));
    InMux I__3092 (
            .O(N__15679),
            .I(N__15659));
    InMux I__3091 (
            .O(N__15678),
            .I(N__15659));
    InMux I__3090 (
            .O(N__15675),
            .I(N__15659));
    Span4Mux_h I__3089 (
            .O(N__15672),
            .I(N__15653));
    InMux I__3088 (
            .O(N__15671),
            .I(N__15650));
    LocalMux I__3087 (
            .O(N__15668),
            .I(N__15645));
    LocalMux I__3086 (
            .O(N__15659),
            .I(N__15645));
    InMux I__3085 (
            .O(N__15658),
            .I(N__15638));
    InMux I__3084 (
            .O(N__15657),
            .I(N__15638));
    InMux I__3083 (
            .O(N__15656),
            .I(N__15638));
    Sp12to4 I__3082 (
            .O(N__15653),
            .I(N__15633));
    LocalMux I__3081 (
            .O(N__15650),
            .I(N__15633));
    Span4Mux_h I__3080 (
            .O(N__15645),
            .I(N__15630));
    LocalMux I__3079 (
            .O(N__15638),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv12 I__3078 (
            .O(N__15633),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__3077 (
            .O(N__15630),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__3076 (
            .O(N__15623),
            .I(N__15620));
    LocalMux I__3075 (
            .O(N__15620),
            .I(\uu2.bitmap_pmux_sn_N_54_mux ));
    InMux I__3074 (
            .O(N__15617),
            .I(N__15614));
    LocalMux I__3073 (
            .O(N__15614),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    CEMux I__3072 (
            .O(N__15611),
            .I(N__15608));
    LocalMux I__3071 (
            .O(N__15608),
            .I(N__15604));
    CEMux I__3070 (
            .O(N__15607),
            .I(N__15601));
    Sp12to4 I__3069 (
            .O(N__15604),
            .I(N__15598));
    LocalMux I__3068 (
            .O(N__15601),
            .I(\uu2.N_31_0 ));
    Odrv12 I__3067 (
            .O(N__15598),
            .I(\uu2.N_31_0 ));
    InMux I__3066 (
            .O(N__15593),
            .I(N__15590));
    LocalMux I__3065 (
            .O(N__15590),
            .I(\uu2.bitmapZ0Z_90 ));
    InMux I__3064 (
            .O(N__15587),
            .I(N__15584));
    LocalMux I__3063 (
            .O(N__15584),
            .I(N__15581));
    Odrv12 I__3062 (
            .O(N__15581),
            .I(\uu2.mem0.N_36 ));
    CascadeMux I__3061 (
            .O(N__15578),
            .I(\uu2.mem0.N_9_cascade_ ));
    InMux I__3060 (
            .O(N__15575),
            .I(N__15572));
    LocalMux I__3059 (
            .O(N__15572),
            .I(\uu2.bitmap_pmux_26_bm_1 ));
    CascadeMux I__3058 (
            .O(N__15569),
            .I(\uu2.bitmap_RNI31F32Z0Z_34_cascade_ ));
    InMux I__3057 (
            .O(N__15566),
            .I(N__15563));
    LocalMux I__3056 (
            .O(N__15563),
            .I(\uu2.w_addr_displaying_RNIBICU6_0Z0Z_2 ));
    CascadeMux I__3055 (
            .O(N__15560),
            .I(\uu2.N_401_cascade_ ));
    InMux I__3054 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__3053 (
            .O(N__15554),
            .I(\uu2.w_addr_displaying_RNIBICU6Z0Z_2 ));
    InMux I__3052 (
            .O(N__15551),
            .I(N__15548));
    LocalMux I__3051 (
            .O(N__15548),
            .I(N__15545));
    Odrv4 I__3050 (
            .O(N__15545),
            .I(\uu2.bitmapZ0Z_111 ));
    CascadeMux I__3049 (
            .O(N__15542),
            .I(\uu2.N_99_cascade_ ));
    InMux I__3048 (
            .O(N__15539),
            .I(N__15536));
    LocalMux I__3047 (
            .O(N__15536),
            .I(\uu2.bitmap_RNI2Q8F1Z0Z_111 ));
    InMux I__3046 (
            .O(N__15533),
            .I(N__15530));
    LocalMux I__3045 (
            .O(N__15530),
            .I(\uu2.bitmap_pmux_sn_N_15 ));
    CascadeMux I__3044 (
            .O(N__15527),
            .I(N__15524));
    InMux I__3043 (
            .O(N__15524),
            .I(N__15521));
    LocalMux I__3042 (
            .O(N__15521),
            .I(bu_rx_data_fast_5));
    InMux I__3041 (
            .O(N__15518),
            .I(N__15515));
    LocalMux I__3040 (
            .O(N__15515),
            .I(bu_rx_data_fast_3));
    CascadeMux I__3039 (
            .O(N__15512),
            .I(\uu2.mem0.N_98_0_cascade_ ));
    InMux I__3038 (
            .O(N__15509),
            .I(N__15506));
    LocalMux I__3037 (
            .O(N__15506),
            .I(\uu2.mem0.G_11_0_0_a3_0_2 ));
    CascadeMux I__3036 (
            .O(N__15503),
            .I(\uu2.mem0.N_62_cascade_ ));
    CascadeMux I__3035 (
            .O(N__15500),
            .I(\Lab_UT.dictrl.g2_1_0_1_cascade_ ));
    InMux I__3034 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__3033 (
            .O(N__15494),
            .I(\Lab_UT.dictrl.N_7_1_0 ));
    CascadeMux I__3032 (
            .O(N__15491),
            .I(N__15488));
    InMux I__3031 (
            .O(N__15488),
            .I(N__15484));
    InMux I__3030 (
            .O(N__15487),
            .I(N__15481));
    LocalMux I__3029 (
            .O(N__15484),
            .I(N__15478));
    LocalMux I__3028 (
            .O(N__15481),
            .I(bu_rx_data_fast_4));
    Odrv4 I__3027 (
            .O(N__15478),
            .I(bu_rx_data_fast_4));
    CascadeMux I__3026 (
            .O(N__15473),
            .I(\Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ));
    InMux I__3025 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__3024 (
            .O(N__15467),
            .I(\Lab_UT.dictrl.next_state18_1_0 ));
    CascadeMux I__3023 (
            .O(N__15464),
            .I(\Lab_UT.dictrl.g1_0_1_cascade_ ));
    InMux I__3022 (
            .O(N__15461),
            .I(N__15458));
    LocalMux I__3021 (
            .O(N__15458),
            .I(\Lab_UT.dictrl.g2_1 ));
    InMux I__3020 (
            .O(N__15455),
            .I(N__15449));
    InMux I__3019 (
            .O(N__15454),
            .I(N__15446));
    InMux I__3018 (
            .O(N__15453),
            .I(N__15441));
    InMux I__3017 (
            .O(N__15452),
            .I(N__15441));
    LocalMux I__3016 (
            .O(N__15449),
            .I(N__15437));
    LocalMux I__3015 (
            .O(N__15446),
            .I(N__15432));
    LocalMux I__3014 (
            .O(N__15441),
            .I(N__15432));
    InMux I__3013 (
            .O(N__15440),
            .I(N__15429));
    Span4Mux_h I__3012 (
            .O(N__15437),
            .I(N__15426));
    Span4Mux_v I__3011 (
            .O(N__15432),
            .I(N__15421));
    LocalMux I__3010 (
            .O(N__15429),
            .I(N__15421));
    Odrv4 I__3009 (
            .O(N__15426),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3008 (
            .O(N__15421),
            .I(\Lab_UT.LdMones ));
    CascadeMux I__3007 (
            .O(N__15416),
            .I(\Lab_UT.dictrl.g0_1_2_0_cascade_ ));
    CascadeMux I__3006 (
            .O(N__15413),
            .I(\Lab_UT.dictrl.N_29_0_0_cascade_ ));
    InMux I__3005 (
            .O(N__15410),
            .I(N__15407));
    LocalMux I__3004 (
            .O(N__15407),
            .I(\Lab_UT.dictrl.N_30_0 ));
    CascadeMux I__3003 (
            .O(N__15404),
            .I(\Lab_UT.dictrl.N_30_0_cascade_ ));
    InMux I__3002 (
            .O(N__15401),
            .I(N__15395));
    InMux I__3001 (
            .O(N__15400),
            .I(N__15395));
    LocalMux I__3000 (
            .O(N__15395),
            .I(\Lab_UT.dictrl.i6_mux_0 ));
    InMux I__2999 (
            .O(N__15392),
            .I(N__15389));
    LocalMux I__2998 (
            .O(N__15389),
            .I(N__15386));
    Odrv4 I__2997 (
            .O(N__15386),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    CascadeMux I__2996 (
            .O(N__15383),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ));
    CascadeMux I__2995 (
            .O(N__15380),
            .I(\Lab_UT.dictrl.dicLdAMones_0_sx_cascade_ ));
    CascadeMux I__2994 (
            .O(N__15377),
            .I(N__15373));
    InMux I__2993 (
            .O(N__15376),
            .I(N__15368));
    InMux I__2992 (
            .O(N__15373),
            .I(N__15368));
    LocalMux I__2991 (
            .O(N__15368),
            .I(N__15365));
    Odrv4 I__2990 (
            .O(N__15365),
            .I(\Lab_UT.dicLdAMones_1 ));
    CascadeMux I__2989 (
            .O(N__15362),
            .I(N__15359));
    InMux I__2988 (
            .O(N__15359),
            .I(N__15356));
    LocalMux I__2987 (
            .O(N__15356),
            .I(\Lab_UT.dictrl.g0_1_3 ));
    CascadeMux I__2986 (
            .O(N__15353),
            .I(N__15349));
    InMux I__2985 (
            .O(N__15352),
            .I(N__15344));
    InMux I__2984 (
            .O(N__15349),
            .I(N__15344));
    LocalMux I__2983 (
            .O(N__15344),
            .I(N__15341));
    Odrv4 I__2982 (
            .O(N__15341),
            .I(\Lab_UT.dicLdSones_1 ));
    CascadeMux I__2981 (
            .O(N__15338),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_ ));
    CascadeMux I__2980 (
            .O(N__15335),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_ ));
    CascadeMux I__2979 (
            .O(N__15332),
            .I(\Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_ ));
    InMux I__2978 (
            .O(N__15329),
            .I(N__15326));
    LocalMux I__2977 (
            .O(N__15326),
            .I(\Lab_UT.dictrl.g0_0_i_a3_2 ));
    CascadeMux I__2976 (
            .O(N__15323),
            .I(\Lab_UT.dictrl.g3_0_cascade_ ));
    InMux I__2975 (
            .O(N__15320),
            .I(N__15317));
    LocalMux I__2974 (
            .O(N__15317),
            .I(\Lab_UT.dictrl.g0_0_0_a3_2 ));
    CascadeMux I__2973 (
            .O(N__15314),
            .I(\Lab_UT.didp.countrce1.q_5_2_cascade_ ));
    CascadeMux I__2972 (
            .O(N__15311),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    InMux I__2971 (
            .O(N__15308),
            .I(N__15296));
    InMux I__2970 (
            .O(N__15307),
            .I(N__15296));
    InMux I__2969 (
            .O(N__15306),
            .I(N__15296));
    InMux I__2968 (
            .O(N__15305),
            .I(N__15296));
    LocalMux I__2967 (
            .O(N__15296),
            .I(N__15293));
    Odrv4 I__2966 (
            .O(N__15293),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    CascadeMux I__2965 (
            .O(N__15290),
            .I(\Lab_UT.didp.countrce1.q_5_3_cascade_ ));
    CascadeMux I__2964 (
            .O(N__15287),
            .I(N__15284));
    InMux I__2963 (
            .O(N__15284),
            .I(N__15281));
    LocalMux I__2962 (
            .O(N__15281),
            .I(N__15278));
    Odrv4 I__2961 (
            .O(N__15278),
            .I(\Lab_UT.didp.countrce1.q_5_1 ));
    CascadeMux I__2960 (
            .O(N__15275),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_ ));
    CascadeMux I__2959 (
            .O(N__15272),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_ ));
    CascadeMux I__2958 (
            .O(N__15269),
            .I(N__15264));
    CascadeMux I__2957 (
            .O(N__15268),
            .I(N__15260));
    InMux I__2956 (
            .O(N__15267),
            .I(N__15257));
    InMux I__2955 (
            .O(N__15264),
            .I(N__15252));
    InMux I__2954 (
            .O(N__15263),
            .I(N__15252));
    InMux I__2953 (
            .O(N__15260),
            .I(N__15249));
    LocalMux I__2952 (
            .O(N__15257),
            .I(\Lab_UT.LdSones ));
    LocalMux I__2951 (
            .O(N__15252),
            .I(\Lab_UT.LdSones ));
    LocalMux I__2950 (
            .O(N__15249),
            .I(\Lab_UT.LdSones ));
    CascadeMux I__2949 (
            .O(N__15242),
            .I(\Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_ ));
    InMux I__2948 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__2947 (
            .O(N__15236),
            .I(N__15233));
    Odrv4 I__2946 (
            .O(N__15233),
            .I(\Lab_UT.bcd2segment3.segment_0Z0Z_0 ));
    InMux I__2945 (
            .O(N__15230),
            .I(N__15224));
    InMux I__2944 (
            .O(N__15229),
            .I(N__15224));
    LocalMux I__2943 (
            .O(N__15224),
            .I(N__15209));
    InMux I__2942 (
            .O(N__15223),
            .I(N__15206));
    InMux I__2941 (
            .O(N__15222),
            .I(N__15203));
    InMux I__2940 (
            .O(N__15221),
            .I(N__15200));
    InMux I__2939 (
            .O(N__15220),
            .I(N__15195));
    InMux I__2938 (
            .O(N__15219),
            .I(N__15195));
    InMux I__2937 (
            .O(N__15218),
            .I(N__15180));
    InMux I__2936 (
            .O(N__15217),
            .I(N__15180));
    InMux I__2935 (
            .O(N__15216),
            .I(N__15180));
    InMux I__2934 (
            .O(N__15215),
            .I(N__15180));
    InMux I__2933 (
            .O(N__15214),
            .I(N__15180));
    InMux I__2932 (
            .O(N__15213),
            .I(N__15180));
    InMux I__2931 (
            .O(N__15212),
            .I(N__15180));
    Span4Mux_h I__2930 (
            .O(N__15209),
            .I(N__15175));
    LocalMux I__2929 (
            .O(N__15206),
            .I(N__15175));
    LocalMux I__2928 (
            .O(N__15203),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__2927 (
            .O(N__15200),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__2926 (
            .O(N__15195),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__2925 (
            .O(N__15180),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__2924 (
            .O(N__15175),
            .I(\Lab_UT.di_Mones_0 ));
    InMux I__2923 (
            .O(N__15164),
            .I(N__15143));
    InMux I__2922 (
            .O(N__15163),
            .I(N__15143));
    InMux I__2921 (
            .O(N__15162),
            .I(N__15143));
    InMux I__2920 (
            .O(N__15161),
            .I(N__15143));
    InMux I__2919 (
            .O(N__15160),
            .I(N__15143));
    InMux I__2918 (
            .O(N__15159),
            .I(N__15143));
    InMux I__2917 (
            .O(N__15158),
            .I(N__15143));
    LocalMux I__2916 (
            .O(N__15143),
            .I(N__15136));
    InMux I__2915 (
            .O(N__15142),
            .I(N__15131));
    InMux I__2914 (
            .O(N__15141),
            .I(N__15131));
    InMux I__2913 (
            .O(N__15140),
            .I(N__15126));
    InMux I__2912 (
            .O(N__15139),
            .I(N__15126));
    Span4Mux_h I__2911 (
            .O(N__15136),
            .I(N__15123));
    LocalMux I__2910 (
            .O(N__15131),
            .I(\Lab_UT.di_Mones_2 ));
    LocalMux I__2909 (
            .O(N__15126),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__2908 (
            .O(N__15123),
            .I(\Lab_UT.di_Mones_2 ));
    CascadeMux I__2907 (
            .O(N__15116),
            .I(N__15106));
    CascadeMux I__2906 (
            .O(N__15115),
            .I(N__15103));
    CascadeMux I__2905 (
            .O(N__15114),
            .I(N__15100));
    CascadeMux I__2904 (
            .O(N__15113),
            .I(N__15097));
    CascadeMux I__2903 (
            .O(N__15112),
            .I(N__15094));
    CascadeMux I__2902 (
            .O(N__15111),
            .I(N__15091));
    CascadeMux I__2901 (
            .O(N__15110),
            .I(N__15088));
    CascadeMux I__2900 (
            .O(N__15109),
            .I(N__15083));
    InMux I__2899 (
            .O(N__15106),
            .I(N__15076));
    InMux I__2898 (
            .O(N__15103),
            .I(N__15076));
    InMux I__2897 (
            .O(N__15100),
            .I(N__15076));
    InMux I__2896 (
            .O(N__15097),
            .I(N__15067));
    InMux I__2895 (
            .O(N__15094),
            .I(N__15067));
    InMux I__2894 (
            .O(N__15091),
            .I(N__15067));
    InMux I__2893 (
            .O(N__15088),
            .I(N__15067));
    InMux I__2892 (
            .O(N__15087),
            .I(N__15064));
    InMux I__2891 (
            .O(N__15086),
            .I(N__15059));
    InMux I__2890 (
            .O(N__15083),
            .I(N__15059));
    LocalMux I__2889 (
            .O(N__15076),
            .I(N__15054));
    LocalMux I__2888 (
            .O(N__15067),
            .I(N__15054));
    LocalMux I__2887 (
            .O(N__15064),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__2886 (
            .O(N__15059),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__2885 (
            .O(N__15054),
            .I(\Lab_UT.di_Mones_3 ));
    CascadeMux I__2884 (
            .O(N__15047),
            .I(N__15043));
    InMux I__2883 (
            .O(N__15046),
            .I(N__15037));
    InMux I__2882 (
            .O(N__15043),
            .I(N__15037));
    CascadeMux I__2881 (
            .O(N__15042),
            .I(N__15034));
    LocalMux I__2880 (
            .O(N__15037),
            .I(N__15029));
    InMux I__2879 (
            .O(N__15034),
            .I(N__15019));
    InMux I__2878 (
            .O(N__15033),
            .I(N__15016));
    InMux I__2877 (
            .O(N__15032),
            .I(N__15013));
    Span4Mux_h I__2876 (
            .O(N__15029),
            .I(N__15010));
    InMux I__2875 (
            .O(N__15028),
            .I(N__15003));
    InMux I__2874 (
            .O(N__15027),
            .I(N__15003));
    InMux I__2873 (
            .O(N__15026),
            .I(N__15003));
    InMux I__2872 (
            .O(N__15025),
            .I(N__14994));
    InMux I__2871 (
            .O(N__15024),
            .I(N__14994));
    InMux I__2870 (
            .O(N__15023),
            .I(N__14994));
    InMux I__2869 (
            .O(N__15022),
            .I(N__14994));
    LocalMux I__2868 (
            .O(N__15019),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2867 (
            .O(N__15016),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2866 (
            .O(N__15013),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv4 I__2865 (
            .O(N__15010),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2864 (
            .O(N__15003),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__2863 (
            .O(N__14994),
            .I(\Lab_UT.di_Mones_1 ));
    CascadeMux I__2862 (
            .O(N__14981),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ));
    CascadeMux I__2861 (
            .O(N__14978),
            .I(N__14975));
    InMux I__2860 (
            .O(N__14975),
            .I(N__14972));
    LocalMux I__2859 (
            .O(N__14972),
            .I(N__14969));
    Span4Mux_h I__2858 (
            .O(N__14969),
            .I(N__14966));
    Odrv4 I__2857 (
            .O(N__14966),
            .I(\uu2.bitmapZ0Z_296 ));
    CascadeMux I__2856 (
            .O(N__14963),
            .I(\Lab_UT.didp.countrce1.q_5_0_cascade_ ));
    InMux I__2855 (
            .O(N__14960),
            .I(N__14957));
    LocalMux I__2854 (
            .O(N__14957),
            .I(\Lab_UT.three_2 ));
    InMux I__2853 (
            .O(N__14954),
            .I(N__14951));
    LocalMux I__2852 (
            .O(N__14951),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_6 ));
    CascadeMux I__2851 (
            .O(N__14948),
            .I(N__14942));
    CascadeMux I__2850 (
            .O(N__14947),
            .I(N__14938));
    InMux I__2849 (
            .O(N__14946),
            .I(N__14935));
    InMux I__2848 (
            .O(N__14945),
            .I(N__14932));
    InMux I__2847 (
            .O(N__14942),
            .I(N__14929));
    InMux I__2846 (
            .O(N__14941),
            .I(N__14926));
    InMux I__2845 (
            .O(N__14938),
            .I(N__14923));
    LocalMux I__2844 (
            .O(N__14935),
            .I(N__14920));
    LocalMux I__2843 (
            .O(N__14932),
            .I(N__14917));
    LocalMux I__2842 (
            .O(N__14929),
            .I(N__14913));
    LocalMux I__2841 (
            .O(N__14926),
            .I(N__14908));
    LocalMux I__2840 (
            .O(N__14923),
            .I(N__14908));
    Span4Mux_h I__2839 (
            .O(N__14920),
            .I(N__14903));
    Span4Mux_v I__2838 (
            .O(N__14917),
            .I(N__14903));
    InMux I__2837 (
            .O(N__14916),
            .I(N__14900));
    Span4Mux_h I__2836 (
            .O(N__14913),
            .I(N__14897));
    Span4Mux_h I__2835 (
            .O(N__14908),
            .I(N__14894));
    Span4Mux_v I__2834 (
            .O(N__14903),
            .I(N__14891));
    LocalMux I__2833 (
            .O(N__14900),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2832 (
            .O(N__14897),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2831 (
            .O(N__14894),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2830 (
            .O(N__14891),
            .I(o_One_Sec_Pulse));
    InMux I__2829 (
            .O(N__14882),
            .I(N__14878));
    InMux I__2828 (
            .O(N__14881),
            .I(N__14875));
    LocalMux I__2827 (
            .O(N__14878),
            .I(N__14872));
    LocalMux I__2826 (
            .O(N__14875),
            .I(N__14867));
    Span4Mux_v I__2825 (
            .O(N__14872),
            .I(N__14864));
    InMux I__2824 (
            .O(N__14871),
            .I(N__14859));
    InMux I__2823 (
            .O(N__14870),
            .I(N__14859));
    Span12Mux_s10_h I__2822 (
            .O(N__14867),
            .I(N__14856));
    Odrv4 I__2821 (
            .O(N__14864),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__2820 (
            .O(N__14859),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv12 I__2819 (
            .O(N__14856),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__2818 (
            .O(N__14849),
            .I(N__14846));
    LocalMux I__2817 (
            .O(N__14846),
            .I(N__14842));
    InMux I__2816 (
            .O(N__14845),
            .I(N__14839));
    Span4Mux_h I__2815 (
            .O(N__14842),
            .I(N__14836));
    LocalMux I__2814 (
            .O(N__14839),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__2813 (
            .O(N__14836),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__2812 (
            .O(N__14831),
            .I(N__14828));
    LocalMux I__2811 (
            .O(N__14828),
            .I(N__14825));
    Span4Mux_h I__2810 (
            .O(N__14825),
            .I(N__14822));
    Odrv4 I__2809 (
            .O(N__14822),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    CascadeMux I__2808 (
            .O(N__14819),
            .I(\uu2.N_97_cascade_ ));
    InMux I__2807 (
            .O(N__14816),
            .I(N__14810));
    InMux I__2806 (
            .O(N__14815),
            .I(N__14810));
    LocalMux I__2805 (
            .O(N__14810),
            .I(\uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2 ));
    InMux I__2804 (
            .O(N__14807),
            .I(N__14804));
    LocalMux I__2803 (
            .O(N__14804),
            .I(\Lab_UT.dictrl.next_alarmstate_1 ));
    InMux I__2802 (
            .O(N__14801),
            .I(N__14798));
    LocalMux I__2801 (
            .O(N__14798),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    InMux I__2800 (
            .O(N__14795),
            .I(N__14779));
    InMux I__2799 (
            .O(N__14794),
            .I(N__14779));
    InMux I__2798 (
            .O(N__14793),
            .I(N__14779));
    InMux I__2797 (
            .O(N__14792),
            .I(N__14779));
    InMux I__2796 (
            .O(N__14791),
            .I(N__14779));
    CascadeMux I__2795 (
            .O(N__14790),
            .I(N__14776));
    LocalMux I__2794 (
            .O(N__14779),
            .I(N__14771));
    InMux I__2793 (
            .O(N__14776),
            .I(N__14764));
    InMux I__2792 (
            .O(N__14775),
            .I(N__14764));
    InMux I__2791 (
            .O(N__14774),
            .I(N__14764));
    Odrv4 I__2790 (
            .O(N__14771),
            .I(\Lab_UT.dictrl.un1_next_alarmstate21_0 ));
    LocalMux I__2789 (
            .O(N__14764),
            .I(\Lab_UT.dictrl.un1_next_alarmstate21_0 ));
    InMux I__2788 (
            .O(N__14759),
            .I(N__14756));
    LocalMux I__2787 (
            .O(N__14756),
            .I(N__14753));
    Span4Mux_h I__2786 (
            .O(N__14753),
            .I(N__14748));
    InMux I__2785 (
            .O(N__14752),
            .I(N__14745));
    InMux I__2784 (
            .O(N__14751),
            .I(N__14742));
    Odrv4 I__2783 (
            .O(N__14748),
            .I(\Lab_UT.di_AStens_1 ));
    LocalMux I__2782 (
            .O(N__14745),
            .I(\Lab_UT.di_AStens_1 ));
    LocalMux I__2781 (
            .O(N__14742),
            .I(\Lab_UT.di_AStens_1 ));
    CascadeMux I__2780 (
            .O(N__14735),
            .I(N__14732));
    InMux I__2779 (
            .O(N__14732),
            .I(N__14729));
    LocalMux I__2778 (
            .O(N__14729),
            .I(N__14726));
    Odrv12 I__2777 (
            .O(N__14726),
            .I(\Lab_UT.sec1Z0Z_1 ));
    InMux I__2776 (
            .O(N__14723),
            .I(N__14719));
    InMux I__2775 (
            .O(N__14722),
            .I(N__14715));
    LocalMux I__2774 (
            .O(N__14719),
            .I(N__14710));
    IoInMux I__2773 (
            .O(N__14718),
            .I(N__14707));
    LocalMux I__2772 (
            .O(N__14715),
            .I(N__14704));
    InMux I__2771 (
            .O(N__14714),
            .I(N__14699));
    InMux I__2770 (
            .O(N__14713),
            .I(N__14699));
    Span4Mux_s3_v I__2769 (
            .O(N__14710),
            .I(N__14696));
    LocalMux I__2768 (
            .O(N__14707),
            .I(N__14693));
    Span4Mux_h I__2767 (
            .O(N__14704),
            .I(N__14690));
    LocalMux I__2766 (
            .O(N__14699),
            .I(N__14687));
    Span4Mux_h I__2765 (
            .O(N__14696),
            .I(N__14682));
    Span4Mux_s3_h I__2764 (
            .O(N__14693),
            .I(N__14682));
    Odrv4 I__2763 (
            .O(N__14690),
            .I(rst));
    Odrv12 I__2762 (
            .O(N__14687),
            .I(rst));
    Odrv4 I__2761 (
            .O(N__14682),
            .I(rst));
    InMux I__2760 (
            .O(N__14675),
            .I(N__14671));
    InMux I__2759 (
            .O(N__14674),
            .I(N__14668));
    LocalMux I__2758 (
            .O(N__14671),
            .I(N__14665));
    LocalMux I__2757 (
            .O(N__14668),
            .I(N__14662));
    Odrv4 I__2756 (
            .O(N__14665),
            .I(\resetGen.un241_ci ));
    Odrv4 I__2755 (
            .O(N__14662),
            .I(\resetGen.un241_ci ));
    CascadeMux I__2754 (
            .O(N__14657),
            .I(N__14654));
    InMux I__2753 (
            .O(N__14654),
            .I(N__14642));
    InMux I__2752 (
            .O(N__14653),
            .I(N__14642));
    InMux I__2751 (
            .O(N__14652),
            .I(N__14642));
    InMux I__2750 (
            .O(N__14651),
            .I(N__14642));
    LocalMux I__2749 (
            .O(N__14642),
            .I(\resetGen.reset_countZ0Z_0 ));
    CascadeMux I__2748 (
            .O(N__14639),
            .I(N__14635));
    InMux I__2747 (
            .O(N__14638),
            .I(N__14631));
    InMux I__2746 (
            .O(N__14635),
            .I(N__14626));
    InMux I__2745 (
            .O(N__14634),
            .I(N__14626));
    LocalMux I__2744 (
            .O(N__14631),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__2743 (
            .O(N__14626),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__2742 (
            .O(N__14621),
            .I(N__14616));
    InMux I__2741 (
            .O(N__14620),
            .I(N__14613));
    InMux I__2740 (
            .O(N__14619),
            .I(N__14610));
    InMux I__2739 (
            .O(N__14616),
            .I(N__14607));
    LocalMux I__2738 (
            .O(N__14613),
            .I(N__14604));
    LocalMux I__2737 (
            .O(N__14610),
            .I(N__14601));
    LocalMux I__2736 (
            .O(N__14607),
            .I(N__14594));
    Span4Mux_v I__2735 (
            .O(N__14604),
            .I(N__14594));
    Span4Mux_v I__2734 (
            .O(N__14601),
            .I(N__14594));
    Odrv4 I__2733 (
            .O(N__14594),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__2732 (
            .O(N__14591),
            .I(N__14582));
    InMux I__2731 (
            .O(N__14590),
            .I(N__14582));
    InMux I__2730 (
            .O(N__14589),
            .I(N__14582));
    LocalMux I__2729 (
            .O(N__14582),
            .I(N__14576));
    InMux I__2728 (
            .O(N__14581),
            .I(N__14573));
    InMux I__2727 (
            .O(N__14580),
            .I(N__14568));
    InMux I__2726 (
            .O(N__14579),
            .I(N__14568));
    Odrv4 I__2725 (
            .O(N__14576),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__2724 (
            .O(N__14573),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__2723 (
            .O(N__14568),
            .I(\resetGen.reset_countZ0Z_4 ));
    CascadeMux I__2722 (
            .O(N__14561),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__2721 (
            .O(N__14558),
            .I(N__14549));
    InMux I__2720 (
            .O(N__14557),
            .I(N__14549));
    InMux I__2719 (
            .O(N__14556),
            .I(N__14549));
    LocalMux I__2718 (
            .O(N__14549),
            .I(N__14544));
    InMux I__2717 (
            .O(N__14548),
            .I(N__14541));
    InMux I__2716 (
            .O(N__14547),
            .I(N__14538));
    Span4Mux_h I__2715 (
            .O(N__14544),
            .I(N__14535));
    LocalMux I__2714 (
            .O(N__14541),
            .I(N__14530));
    LocalMux I__2713 (
            .O(N__14538),
            .I(N__14530));
    Span4Mux_v I__2712 (
            .O(N__14535),
            .I(N__14527));
    Span4Mux_v I__2711 (
            .O(N__14530),
            .I(N__14524));
    Odrv4 I__2710 (
            .O(N__14527),
            .I(\resetGen.escKeyZ0 ));
    Odrv4 I__2709 (
            .O(N__14524),
            .I(\resetGen.escKeyZ0 ));
    InMux I__2708 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__2707 (
            .O(N__14516),
            .I(N__14513));
    Span4Mux_v I__2706 (
            .O(N__14513),
            .I(N__14509));
    InMux I__2705 (
            .O(N__14512),
            .I(N__14506));
    Span4Mux_h I__2704 (
            .O(N__14509),
            .I(N__14503));
    LocalMux I__2703 (
            .O(N__14506),
            .I(\resetGen.reset_countZ0Z_3 ));
    Odrv4 I__2702 (
            .O(N__14503),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__2701 (
            .O(N__14498),
            .I(N__14493));
    InMux I__2700 (
            .O(N__14497),
            .I(N__14489));
    InMux I__2699 (
            .O(N__14496),
            .I(N__14484));
    InMux I__2698 (
            .O(N__14493),
            .I(N__14484));
    InMux I__2697 (
            .O(N__14492),
            .I(N__14480));
    LocalMux I__2696 (
            .O(N__14489),
            .I(N__14475));
    LocalMux I__2695 (
            .O(N__14484),
            .I(N__14475));
    InMux I__2694 (
            .O(N__14483),
            .I(N__14472));
    LocalMux I__2693 (
            .O(N__14480),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__2692 (
            .O(N__14475),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__2691 (
            .O(N__14472),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__2690 (
            .O(N__14465),
            .I(N__14461));
    CascadeMux I__2689 (
            .O(N__14464),
            .I(N__14456));
    InMux I__2688 (
            .O(N__14461),
            .I(N__14451));
    InMux I__2687 (
            .O(N__14460),
            .I(N__14451));
    InMux I__2686 (
            .O(N__14459),
            .I(N__14446));
    InMux I__2685 (
            .O(N__14456),
            .I(N__14446));
    LocalMux I__2684 (
            .O(N__14451),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__2683 (
            .O(N__14446),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__2682 (
            .O(N__14441),
            .I(N__14438));
    LocalMux I__2681 (
            .O(N__14438),
            .I(\uu2.vbuf_w_addr_user.un448_ci_0 ));
    InMux I__2680 (
            .O(N__14435),
            .I(N__14432));
    LocalMux I__2679 (
            .O(N__14432),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__2678 (
            .O(N__14429),
            .I(N__14426));
    InMux I__2677 (
            .O(N__14426),
            .I(N__14423));
    LocalMux I__2676 (
            .O(N__14423),
            .I(\Lab_UT.bcd2segment2.segment_0Z0Z_0 ));
    CascadeMux I__2675 (
            .O(N__14420),
            .I(N__14417));
    InMux I__2674 (
            .O(N__14417),
            .I(N__14414));
    LocalMux I__2673 (
            .O(N__14414),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    InMux I__2672 (
            .O(N__14411),
            .I(N__14405));
    InMux I__2671 (
            .O(N__14410),
            .I(N__14405));
    LocalMux I__2670 (
            .O(N__14405),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    CascadeMux I__2669 (
            .O(N__14402),
            .I(\uu2.bitmap_pmux_sn_N_11_cascade_ ));
    InMux I__2668 (
            .O(N__14399),
            .I(N__14396));
    LocalMux I__2667 (
            .O(N__14396),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__2666 (
            .O(N__14393),
            .I(N__14390));
    LocalMux I__2665 (
            .O(N__14390),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__2664 (
            .O(N__14387),
            .I(N__14381));
    InMux I__2663 (
            .O(N__14386),
            .I(N__14374));
    InMux I__2662 (
            .O(N__14385),
            .I(N__14374));
    InMux I__2661 (
            .O(N__14384),
            .I(N__14374));
    LocalMux I__2660 (
            .O(N__14381),
            .I(N__14371));
    LocalMux I__2659 (
            .O(N__14374),
            .I(N__14363));
    Span4Mux_v I__2658 (
            .O(N__14371),
            .I(N__14363));
    InMux I__2657 (
            .O(N__14370),
            .I(N__14360));
    InMux I__2656 (
            .O(N__14369),
            .I(N__14355));
    InMux I__2655 (
            .O(N__14368),
            .I(N__14355));
    Odrv4 I__2654 (
            .O(N__14363),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__2653 (
            .O(N__14360),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__2652 (
            .O(N__14355),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__2651 (
            .O(N__14348),
            .I(N__14345));
    InMux I__2650 (
            .O(N__14345),
            .I(N__14342));
    LocalMux I__2649 (
            .O(N__14342),
            .I(N__14336));
    CascadeMux I__2648 (
            .O(N__14341),
            .I(N__14333));
    InMux I__2647 (
            .O(N__14340),
            .I(N__14329));
    InMux I__2646 (
            .O(N__14339),
            .I(N__14326));
    Span4Mux_h I__2645 (
            .O(N__14336),
            .I(N__14323));
    InMux I__2644 (
            .O(N__14333),
            .I(N__14320));
    InMux I__2643 (
            .O(N__14332),
            .I(N__14317));
    LocalMux I__2642 (
            .O(N__14329),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__2641 (
            .O(N__14326),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__2640 (
            .O(N__14323),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__2639 (
            .O(N__14320),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__2638 (
            .O(N__14317),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__2637 (
            .O(N__14306),
            .I(N__14302));
    InMux I__2636 (
            .O(N__14305),
            .I(N__14298));
    InMux I__2635 (
            .O(N__14302),
            .I(N__14295));
    CascadeMux I__2634 (
            .O(N__14301),
            .I(N__14291));
    LocalMux I__2633 (
            .O(N__14298),
            .I(N__14287));
    LocalMux I__2632 (
            .O(N__14295),
            .I(N__14284));
    InMux I__2631 (
            .O(N__14294),
            .I(N__14280));
    InMux I__2630 (
            .O(N__14291),
            .I(N__14275));
    InMux I__2629 (
            .O(N__14290),
            .I(N__14275));
    Span4Mux_v I__2628 (
            .O(N__14287),
            .I(N__14272));
    Span4Mux_h I__2627 (
            .O(N__14284),
            .I(N__14269));
    InMux I__2626 (
            .O(N__14283),
            .I(N__14266));
    LocalMux I__2625 (
            .O(N__14280),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__2624 (
            .O(N__14275),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__2623 (
            .O(N__14272),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__2622 (
            .O(N__14269),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__2621 (
            .O(N__14266),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__2620 (
            .O(N__14255),
            .I(N__14252));
    InMux I__2619 (
            .O(N__14252),
            .I(N__14249));
    LocalMux I__2618 (
            .O(N__14249),
            .I(N__14245));
    InMux I__2617 (
            .O(N__14248),
            .I(N__14241));
    Span4Mux_h I__2616 (
            .O(N__14245),
            .I(N__14238));
    CascadeMux I__2615 (
            .O(N__14244),
            .I(N__14235));
    LocalMux I__2614 (
            .O(N__14241),
            .I(N__14231));
    Sp12to4 I__2613 (
            .O(N__14238),
            .I(N__14228));
    InMux I__2612 (
            .O(N__14235),
            .I(N__14223));
    InMux I__2611 (
            .O(N__14234),
            .I(N__14223));
    Odrv4 I__2610 (
            .O(N__14231),
            .I(\uu2.w_addr_userZ0Z_3 ));
    Odrv12 I__2609 (
            .O(N__14228),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__2608 (
            .O(N__14223),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__2607 (
            .O(N__14216),
            .I(N__14213));
    InMux I__2606 (
            .O(N__14213),
            .I(N__14210));
    LocalMux I__2605 (
            .O(N__14210),
            .I(N__14204));
    InMux I__2604 (
            .O(N__14209),
            .I(N__14199));
    InMux I__2603 (
            .O(N__14208),
            .I(N__14199));
    InMux I__2602 (
            .O(N__14207),
            .I(N__14196));
    Span4Mux_h I__2601 (
            .O(N__14204),
            .I(N__14191));
    LocalMux I__2600 (
            .O(N__14199),
            .I(N__14191));
    LocalMux I__2599 (
            .O(N__14196),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__2598 (
            .O(N__14191),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__2597 (
            .O(N__14186),
            .I(N__14183));
    InMux I__2596 (
            .O(N__14183),
            .I(N__14178));
    CascadeMux I__2595 (
            .O(N__14182),
            .I(N__14174));
    InMux I__2594 (
            .O(N__14181),
            .I(N__14170));
    LocalMux I__2593 (
            .O(N__14178),
            .I(N__14167));
    CascadeMux I__2592 (
            .O(N__14177),
            .I(N__14164));
    InMux I__2591 (
            .O(N__14174),
            .I(N__14159));
    InMux I__2590 (
            .O(N__14173),
            .I(N__14159));
    LocalMux I__2589 (
            .O(N__14170),
            .I(N__14154));
    Span4Mux_h I__2588 (
            .O(N__14167),
            .I(N__14154));
    InMux I__2587 (
            .O(N__14164),
            .I(N__14151));
    LocalMux I__2586 (
            .O(N__14159),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__2585 (
            .O(N__14154),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__2584 (
            .O(N__14151),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__2583 (
            .O(N__14144),
            .I(\uu2.un426_ci_3_cascade_ ));
    CascadeMux I__2582 (
            .O(N__14141),
            .I(N__14138));
    InMux I__2581 (
            .O(N__14138),
            .I(N__14135));
    LocalMux I__2580 (
            .O(N__14135),
            .I(N__14131));
    InMux I__2579 (
            .O(N__14134),
            .I(N__14128));
    Odrv4 I__2578 (
            .O(N__14131),
            .I(\uu2.un426_ci_3 ));
    LocalMux I__2577 (
            .O(N__14128),
            .I(\uu2.un426_ci_3 ));
    InMux I__2576 (
            .O(N__14123),
            .I(N__14112));
    InMux I__2575 (
            .O(N__14122),
            .I(N__14112));
    InMux I__2574 (
            .O(N__14121),
            .I(N__14112));
    InMux I__2573 (
            .O(N__14120),
            .I(N__14107));
    InMux I__2572 (
            .O(N__14119),
            .I(N__14107));
    LocalMux I__2571 (
            .O(N__14112),
            .I(N__14104));
    LocalMux I__2570 (
            .O(N__14107),
            .I(N__14101));
    Span4Mux_h I__2569 (
            .O(N__14104),
            .I(N__14098));
    Span4Mux_h I__2568 (
            .O(N__14101),
            .I(N__14095));
    Odrv4 I__2567 (
            .O(N__14098),
            .I(\uu2.un404_ci ));
    Odrv4 I__2566 (
            .O(N__14095),
            .I(\uu2.un404_ci ));
    CascadeMux I__2565 (
            .O(N__14090),
            .I(N__14087));
    InMux I__2564 (
            .O(N__14087),
            .I(N__14082));
    InMux I__2563 (
            .O(N__14086),
            .I(N__14079));
    InMux I__2562 (
            .O(N__14085),
            .I(N__14076));
    LocalMux I__2561 (
            .O(N__14082),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__2560 (
            .O(N__14079),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__2559 (
            .O(N__14076),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CEMux I__2558 (
            .O(N__14069),
            .I(N__14066));
    LocalMux I__2557 (
            .O(N__14066),
            .I(N__14063));
    Span4Mux_v I__2556 (
            .O(N__14063),
            .I(N__14060));
    Span4Mux_s0_v I__2555 (
            .O(N__14060),
            .I(N__14057));
    Odrv4 I__2554 (
            .O(N__14057),
            .I(\uu2.un28_w_addr_user_i_0 ));
    SRMux I__2553 (
            .O(N__14054),
            .I(N__14051));
    LocalMux I__2552 (
            .O(N__14051),
            .I(N__14048));
    Span4Mux_s1_v I__2551 (
            .O(N__14048),
            .I(N__14043));
    SRMux I__2550 (
            .O(N__14047),
            .I(N__14040));
    SRMux I__2549 (
            .O(N__14046),
            .I(N__14037));
    Span4Mux_h I__2548 (
            .O(N__14043),
            .I(N__14032));
    LocalMux I__2547 (
            .O(N__14040),
            .I(N__14032));
    LocalMux I__2546 (
            .O(N__14037),
            .I(N__14029));
    Span4Mux_h I__2545 (
            .O(N__14032),
            .I(N__14026));
    Odrv12 I__2544 (
            .O(N__14029),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    Odrv4 I__2543 (
            .O(N__14026),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    CascadeMux I__2542 (
            .O(N__14021),
            .I(N__14018));
    InMux I__2541 (
            .O(N__14018),
            .I(N__14015));
    LocalMux I__2540 (
            .O(N__14015),
            .I(N__14012));
    Span4Mux_s3_v I__2539 (
            .O(N__14012),
            .I(N__14009));
    Span4Mux_h I__2538 (
            .O(N__14009),
            .I(N__14006));
    Odrv4 I__2537 (
            .O(N__14006),
            .I(\uu2.mem0.w_addr_6 ));
    CascadeMux I__2536 (
            .O(N__14003),
            .I(N__14000));
    InMux I__2535 (
            .O(N__14000),
            .I(N__13997));
    LocalMux I__2534 (
            .O(N__13997),
            .I(N__13994));
    Span4Mux_h I__2533 (
            .O(N__13994),
            .I(N__13991));
    Odrv4 I__2532 (
            .O(N__13991),
            .I(\uu2.mem0.w_addr_7 ));
    InMux I__2531 (
            .O(N__13988),
            .I(N__13985));
    LocalMux I__2530 (
            .O(N__13985),
            .I(\uu2.mem0.bitmap_pmux_sn_N_42 ));
    InMux I__2529 (
            .O(N__13982),
            .I(N__13979));
    LocalMux I__2528 (
            .O(N__13979),
            .I(N__13976));
    Odrv4 I__2527 (
            .O(N__13976),
            .I(\uu2.un1_w_user_lf_0_0 ));
    CascadeMux I__2526 (
            .O(N__13973),
            .I(N__13970));
    InMux I__2525 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__2524 (
            .O(N__13967),
            .I(N__13964));
    Span4Mux_s1_v I__2523 (
            .O(N__13964),
            .I(N__13961));
    Span4Mux_v I__2522 (
            .O(N__13961),
            .I(N__13958));
    Odrv4 I__2521 (
            .O(N__13958),
            .I(\uu2.un1_w_user_lfZ0Z_4 ));
    InMux I__2520 (
            .O(N__13955),
            .I(N__13952));
    LocalMux I__2519 (
            .O(N__13952),
            .I(\uu2.un20_w_addr_userZ0Z_1 ));
    InMux I__2518 (
            .O(N__13949),
            .I(N__13943));
    InMux I__2517 (
            .O(N__13948),
            .I(N__13943));
    LocalMux I__2516 (
            .O(N__13943),
            .I(\uu2.un3_w_addr_user ));
    CascadeMux I__2515 (
            .O(N__13940),
            .I(\uu2.un20_w_addr_userZ0Z_1_cascade_ ));
    CascadeMux I__2514 (
            .O(N__13937),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2_cascade_ ));
    InMux I__2513 (
            .O(N__13934),
            .I(N__13921));
    InMux I__2512 (
            .O(N__13933),
            .I(N__13921));
    InMux I__2511 (
            .O(N__13932),
            .I(N__13921));
    InMux I__2510 (
            .O(N__13931),
            .I(N__13912));
    InMux I__2509 (
            .O(N__13930),
            .I(N__13912));
    InMux I__2508 (
            .O(N__13929),
            .I(N__13912));
    InMux I__2507 (
            .O(N__13928),
            .I(N__13912));
    LocalMux I__2506 (
            .O(N__13921),
            .I(\uu2.un28_w_addr_user_i ));
    LocalMux I__2505 (
            .O(N__13912),
            .I(\uu2.un28_w_addr_user_i ));
    InMux I__2504 (
            .O(N__13907),
            .I(N__13904));
    LocalMux I__2503 (
            .O(N__13904),
            .I(N__13901));
    Odrv4 I__2502 (
            .O(N__13901),
            .I(\uu2.un3_w_addr_user_5 ));
    InMux I__2501 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__2500 (
            .O(N__13895),
            .I(N__13892));
    Span4Mux_v I__2499 (
            .O(N__13892),
            .I(N__13889));
    Odrv4 I__2498 (
            .O(N__13889),
            .I(bu_rx_data_fast_6));
    CascadeMux I__2497 (
            .O(N__13886),
            .I(N__13883));
    InMux I__2496 (
            .O(N__13883),
            .I(N__13880));
    LocalMux I__2495 (
            .O(N__13880),
            .I(bu_rx_data_fast_7));
    InMux I__2494 (
            .O(N__13877),
            .I(N__13868));
    InMux I__2493 (
            .O(N__13876),
            .I(N__13868));
    InMux I__2492 (
            .O(N__13875),
            .I(N__13868));
    LocalMux I__2491 (
            .O(N__13868),
            .I(N__13864));
    InMux I__2490 (
            .O(N__13867),
            .I(N__13861));
    Span4Mux_s3_v I__2489 (
            .O(N__13864),
            .I(N__13856));
    LocalMux I__2488 (
            .O(N__13861),
            .I(N__13856));
    Odrv4 I__2487 (
            .O(N__13856),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__2486 (
            .O(N__13853),
            .I(N__13850));
    LocalMux I__2485 (
            .O(N__13850),
            .I(\Lab_UT.dictrl.g2_1_0_0 ));
    InMux I__2484 (
            .O(N__13847),
            .I(N__13837));
    InMux I__2483 (
            .O(N__13846),
            .I(N__13837));
    InMux I__2482 (
            .O(N__13845),
            .I(N__13828));
    InMux I__2481 (
            .O(N__13844),
            .I(N__13828));
    InMux I__2480 (
            .O(N__13843),
            .I(N__13828));
    InMux I__2479 (
            .O(N__13842),
            .I(N__13828));
    LocalMux I__2478 (
            .O(N__13837),
            .I(N__13823));
    LocalMux I__2477 (
            .O(N__13828),
            .I(N__13823));
    Odrv4 I__2476 (
            .O(N__13823),
            .I(\Lab_UT.nine ));
    CascadeMux I__2475 (
            .O(N__13820),
            .I(N__13814));
    InMux I__2474 (
            .O(N__13819),
            .I(N__13809));
    InMux I__2473 (
            .O(N__13818),
            .I(N__13809));
    InMux I__2472 (
            .O(N__13817),
            .I(N__13806));
    InMux I__2471 (
            .O(N__13814),
            .I(N__13803));
    LocalMux I__2470 (
            .O(N__13809),
            .I(N__13796));
    LocalMux I__2469 (
            .O(N__13806),
            .I(N__13796));
    LocalMux I__2468 (
            .O(N__13803),
            .I(N__13796));
    Odrv4 I__2467 (
            .O(N__13796),
            .I(\Lab_UT.five ));
    CascadeMux I__2466 (
            .O(N__13793),
            .I(N__13787));
    InMux I__2465 (
            .O(N__13792),
            .I(N__13777));
    InMux I__2464 (
            .O(N__13791),
            .I(N__13777));
    InMux I__2463 (
            .O(N__13790),
            .I(N__13777));
    InMux I__2462 (
            .O(N__13787),
            .I(N__13777));
    CascadeMux I__2461 (
            .O(N__13786),
            .I(N__13773));
    LocalMux I__2460 (
            .O(N__13777),
            .I(N__13770));
    InMux I__2459 (
            .O(N__13776),
            .I(N__13765));
    InMux I__2458 (
            .O(N__13773),
            .I(N__13765));
    Span4Mux_h I__2457 (
            .O(N__13770),
            .I(N__13759));
    LocalMux I__2456 (
            .O(N__13765),
            .I(N__13759));
    InMux I__2455 (
            .O(N__13764),
            .I(N__13756));
    Span4Mux_v I__2454 (
            .O(N__13759),
            .I(N__13753));
    LocalMux I__2453 (
            .O(N__13756),
            .I(N__13750));
    Span4Mux_h I__2452 (
            .O(N__13753),
            .I(N__13747));
    Span4Mux_v I__2451 (
            .O(N__13750),
            .I(N__13744));
    Odrv4 I__2450 (
            .O(N__13747),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    Odrv4 I__2449 (
            .O(N__13744),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    InMux I__2448 (
            .O(N__13739),
            .I(N__13734));
    InMux I__2447 (
            .O(N__13738),
            .I(N__13729));
    InMux I__2446 (
            .O(N__13737),
            .I(N__13729));
    LocalMux I__2445 (
            .O(N__13734),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__2444 (
            .O(N__13729),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__2443 (
            .O(N__13724),
            .I(N__13719));
    InMux I__2442 (
            .O(N__13723),
            .I(N__13714));
    InMux I__2441 (
            .O(N__13722),
            .I(N__13714));
    InMux I__2440 (
            .O(N__13719),
            .I(N__13710));
    LocalMux I__2439 (
            .O(N__13714),
            .I(N__13707));
    InMux I__2438 (
            .O(N__13713),
            .I(N__13704));
    LocalMux I__2437 (
            .O(N__13710),
            .I(N__13701));
    Span4Mux_v I__2436 (
            .O(N__13707),
            .I(N__13698));
    LocalMux I__2435 (
            .O(N__13704),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    Odrv12 I__2434 (
            .O(N__13701),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    Odrv4 I__2433 (
            .O(N__13698),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__2432 (
            .O(N__13691),
            .I(N__13686));
    InMux I__2431 (
            .O(N__13690),
            .I(N__13681));
    InMux I__2430 (
            .O(N__13689),
            .I(N__13681));
    LocalMux I__2429 (
            .O(N__13686),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__2428 (
            .O(N__13681),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__2427 (
            .O(N__13676),
            .I(N__13673));
    LocalMux I__2426 (
            .O(N__13673),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__2425 (
            .O(N__13670),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__2424 (
            .O(N__13667),
            .I(N__13663));
    InMux I__2423 (
            .O(N__13666),
            .I(N__13660));
    LocalMux I__2422 (
            .O(N__13663),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__2421 (
            .O(N__13660),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__2420 (
            .O(N__13655),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__2419 (
            .O(N__13652),
            .I(N__13647));
    InMux I__2418 (
            .O(N__13651),
            .I(N__13642));
    InMux I__2417 (
            .O(N__13650),
            .I(N__13642));
    LocalMux I__2416 (
            .O(N__13647),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__2415 (
            .O(N__13642),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__2414 (
            .O(N__13637),
            .I(N__13634));
    LocalMux I__2413 (
            .O(N__13634),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__2412 (
            .O(N__13631),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__2411 (
            .O(N__13628),
            .I(N__13624));
    CascadeMux I__2410 (
            .O(N__13627),
            .I(N__13620));
    LocalMux I__2409 (
            .O(N__13624),
            .I(N__13616));
    InMux I__2408 (
            .O(N__13623),
            .I(N__13613));
    InMux I__2407 (
            .O(N__13620),
            .I(N__13608));
    InMux I__2406 (
            .O(N__13619),
            .I(N__13608));
    Odrv4 I__2405 (
            .O(N__13616),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__2404 (
            .O(N__13613),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__2403 (
            .O(N__13608),
            .I(\buart.Z_rx.ser_clk ));
    InMux I__2402 (
            .O(N__13601),
            .I(N__13595));
    InMux I__2401 (
            .O(N__13600),
            .I(N__13590));
    InMux I__2400 (
            .O(N__13599),
            .I(N__13590));
    CascadeMux I__2399 (
            .O(N__13598),
            .I(N__13582));
    LocalMux I__2398 (
            .O(N__13595),
            .I(N__13577));
    LocalMux I__2397 (
            .O(N__13590),
            .I(N__13574));
    InMux I__2396 (
            .O(N__13589),
            .I(N__13571));
    InMux I__2395 (
            .O(N__13588),
            .I(N__13568));
    InMux I__2394 (
            .O(N__13587),
            .I(N__13565));
    InMux I__2393 (
            .O(N__13586),
            .I(N__13560));
    InMux I__2392 (
            .O(N__13585),
            .I(N__13560));
    InMux I__2391 (
            .O(N__13582),
            .I(N__13553));
    InMux I__2390 (
            .O(N__13581),
            .I(N__13553));
    InMux I__2389 (
            .O(N__13580),
            .I(N__13553));
    Span4Mux_v I__2388 (
            .O(N__13577),
            .I(N__13550));
    Span4Mux_v I__2387 (
            .O(N__13574),
            .I(N__13547));
    LocalMux I__2386 (
            .O(N__13571),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2385 (
            .O(N__13568),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2384 (
            .O(N__13565),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2383 (
            .O(N__13560),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2382 (
            .O(N__13553),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__2381 (
            .O(N__13550),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__2380 (
            .O(N__13547),
            .I(\buart.Z_rx.startbit ));
    InMux I__2379 (
            .O(N__13532),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__2378 (
            .O(N__13529),
            .I(N__13525));
    CascadeMux I__2377 (
            .O(N__13528),
            .I(N__13522));
    InMux I__2376 (
            .O(N__13525),
            .I(N__13519));
    InMux I__2375 (
            .O(N__13522),
            .I(N__13516));
    LocalMux I__2374 (
            .O(N__13519),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__2373 (
            .O(N__13516),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__2372 (
            .O(N__13511),
            .I(\Lab_UT.dictrl.g2_0_1_0_cascade_ ));
    InMux I__2371 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__2370 (
            .O(N__13505),
            .I(\Lab_UT.didp.countrce4.q_5_0 ));
    InMux I__2369 (
            .O(N__13502),
            .I(N__13499));
    LocalMux I__2368 (
            .O(N__13499),
            .I(N__13494));
    InMux I__2367 (
            .O(N__13498),
            .I(N__13491));
    InMux I__2366 (
            .O(N__13497),
            .I(N__13488));
    Span4Mux_v I__2365 (
            .O(N__13494),
            .I(N__13485));
    LocalMux I__2364 (
            .O(N__13491),
            .I(uu0_sec_clkD));
    LocalMux I__2363 (
            .O(N__13488),
            .I(uu0_sec_clkD));
    Odrv4 I__2362 (
            .O(N__13485),
            .I(uu0_sec_clkD));
    CEMux I__2361 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__2360 (
            .O(N__13475),
            .I(N__13472));
    Sp12to4 I__2359 (
            .O(N__13472),
            .I(N__13469));
    Odrv12 I__2358 (
            .O(N__13469),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    InMux I__2357 (
            .O(N__13466),
            .I(N__13460));
    InMux I__2356 (
            .O(N__13465),
            .I(N__13460));
    LocalMux I__2355 (
            .O(N__13460),
            .I(\Lab_UT.didp.ce_11_0_2 ));
    CascadeMux I__2354 (
            .O(N__13457),
            .I(\Lab_UT.didp.un26_ce_0_cascade_ ));
    InMux I__2353 (
            .O(N__13454),
            .I(N__13443));
    InMux I__2352 (
            .O(N__13453),
            .I(N__13443));
    InMux I__2351 (
            .O(N__13452),
            .I(N__13438));
    InMux I__2350 (
            .O(N__13451),
            .I(N__13438));
    InMux I__2349 (
            .O(N__13450),
            .I(N__13433));
    InMux I__2348 (
            .O(N__13449),
            .I(N__13433));
    InMux I__2347 (
            .O(N__13448),
            .I(N__13430));
    LocalMux I__2346 (
            .O(N__13443),
            .I(N__13427));
    LocalMux I__2345 (
            .O(N__13438),
            .I(N__13422));
    LocalMux I__2344 (
            .O(N__13433),
            .I(N__13422));
    LocalMux I__2343 (
            .O(N__13430),
            .I(N__13419));
    Span12Mux_s5_h I__2342 (
            .O(N__13427),
            .I(N__13416));
    Span4Mux_v I__2341 (
            .O(N__13422),
            .I(N__13413));
    Odrv4 I__2340 (
            .O(N__13419),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    Odrv12 I__2339 (
            .O(N__13416),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    Odrv4 I__2338 (
            .O(N__13413),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    CascadeMux I__2337 (
            .O(N__13406),
            .I(\Lab_UT.didp.ce_12_0_3_cascade_ ));
    InMux I__2336 (
            .O(N__13403),
            .I(N__13400));
    LocalMux I__2335 (
            .O(N__13400),
            .I(\Lab_UT.didp.un26_ce_0 ));
    InMux I__2334 (
            .O(N__13397),
            .I(N__13391));
    InMux I__2333 (
            .O(N__13396),
            .I(N__13391));
    LocalMux I__2332 (
            .O(N__13391),
            .I(N__13384));
    InMux I__2331 (
            .O(N__13390),
            .I(N__13375));
    InMux I__2330 (
            .O(N__13389),
            .I(N__13375));
    InMux I__2329 (
            .O(N__13388),
            .I(N__13375));
    InMux I__2328 (
            .O(N__13387),
            .I(N__13375));
    Span4Mux_h I__2327 (
            .O(N__13384),
            .I(N__13372));
    LocalMux I__2326 (
            .O(N__13375),
            .I(N__13369));
    Odrv4 I__2325 (
            .O(N__13372),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv4 I__2324 (
            .O(N__13369),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    CascadeMux I__2323 (
            .O(N__13364),
            .I(N__13361));
    InMux I__2322 (
            .O(N__13361),
            .I(N__13354));
    InMux I__2321 (
            .O(N__13360),
            .I(N__13354));
    InMux I__2320 (
            .O(N__13359),
            .I(N__13351));
    LocalMux I__2319 (
            .O(N__13354),
            .I(N__13348));
    LocalMux I__2318 (
            .O(N__13351),
            .I(N__13343));
    Span4Mux_h I__2317 (
            .O(N__13348),
            .I(N__13343));
    Odrv4 I__2316 (
            .O(N__13343),
            .I(\Lab_UT.nine_0 ));
    CascadeMux I__2315 (
            .O(N__13340),
            .I(N__13336));
    InMux I__2314 (
            .O(N__13339),
            .I(N__13329));
    InMux I__2313 (
            .O(N__13336),
            .I(N__13329));
    CascadeMux I__2312 (
            .O(N__13335),
            .I(N__13323));
    CascadeMux I__2311 (
            .O(N__13334),
            .I(N__13320));
    LocalMux I__2310 (
            .O(N__13329),
            .I(N__13317));
    InMux I__2309 (
            .O(N__13328),
            .I(N__13312));
    InMux I__2308 (
            .O(N__13327),
            .I(N__13312));
    InMux I__2307 (
            .O(N__13326),
            .I(N__13309));
    InMux I__2306 (
            .O(N__13323),
            .I(N__13306));
    InMux I__2305 (
            .O(N__13320),
            .I(N__13303));
    Span4Mux_h I__2304 (
            .O(N__13317),
            .I(N__13300));
    LocalMux I__2303 (
            .O(N__13312),
            .I(N__13297));
    LocalMux I__2302 (
            .O(N__13309),
            .I(N__13290));
    LocalMux I__2301 (
            .O(N__13306),
            .I(N__13290));
    LocalMux I__2300 (
            .O(N__13303),
            .I(N__13290));
    Odrv4 I__2299 (
            .O(N__13300),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    Odrv4 I__2298 (
            .O(N__13297),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    Odrv12 I__2297 (
            .O(N__13290),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    CascadeMux I__2296 (
            .O(N__13283),
            .I(N__13280));
    InMux I__2295 (
            .O(N__13280),
            .I(N__13265));
    InMux I__2294 (
            .O(N__13279),
            .I(N__13265));
    InMux I__2293 (
            .O(N__13278),
            .I(N__13265));
    InMux I__2292 (
            .O(N__13277),
            .I(N__13265));
    InMux I__2291 (
            .O(N__13276),
            .I(N__13262));
    InMux I__2290 (
            .O(N__13275),
            .I(N__13257));
    InMux I__2289 (
            .O(N__13274),
            .I(N__13257));
    LocalMux I__2288 (
            .O(N__13265),
            .I(N__13254));
    LocalMux I__2287 (
            .O(N__13262),
            .I(N__13249));
    LocalMux I__2286 (
            .O(N__13257),
            .I(N__13249));
    Sp12to4 I__2285 (
            .O(N__13254),
            .I(N__13246));
    Span4Mux_h I__2284 (
            .O(N__13249),
            .I(N__13243));
    Odrv12 I__2283 (
            .O(N__13246),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    Odrv4 I__2282 (
            .O(N__13243),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    CascadeMux I__2281 (
            .O(N__13238),
            .I(\Lab_UT.three_2_2_cascade_ ));
    CascadeMux I__2280 (
            .O(N__13235),
            .I(\Lab_UT.didp.countrce4.q_5_2_cascade_ ));
    CascadeMux I__2279 (
            .O(N__13232),
            .I(\Lab_UT.didp.reset_12_3_3_cascade_ ));
    CascadeMux I__2278 (
            .O(N__13229),
            .I(\Lab_UT.didp.reset_12_1_3_cascade_ ));
    CascadeMux I__2277 (
            .O(N__13226),
            .I(N__13222));
    CascadeMux I__2276 (
            .O(N__13225),
            .I(N__13217));
    InMux I__2275 (
            .O(N__13222),
            .I(N__13210));
    InMux I__2274 (
            .O(N__13221),
            .I(N__13210));
    InMux I__2273 (
            .O(N__13220),
            .I(N__13201));
    InMux I__2272 (
            .O(N__13217),
            .I(N__13201));
    InMux I__2271 (
            .O(N__13216),
            .I(N__13201));
    InMux I__2270 (
            .O(N__13215),
            .I(N__13201));
    LocalMux I__2269 (
            .O(N__13210),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    LocalMux I__2268 (
            .O(N__13201),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    CascadeMux I__2267 (
            .O(N__13196),
            .I(\Lab_UT.didp.countrce4.un20_qPone_cascade_ ));
    InMux I__2266 (
            .O(N__13193),
            .I(N__13189));
    InMux I__2265 (
            .O(N__13192),
            .I(N__13186));
    LocalMux I__2264 (
            .O(N__13189),
            .I(\Lab_UT.didp.countrce4.q_5_3 ));
    LocalMux I__2263 (
            .O(N__13186),
            .I(\Lab_UT.didp.countrce4.q_5_3 ));
    CascadeMux I__2262 (
            .O(N__13181),
            .I(N__13177));
    InMux I__2261 (
            .O(N__13180),
            .I(N__13174));
    InMux I__2260 (
            .O(N__13177),
            .I(N__13171));
    LocalMux I__2259 (
            .O(N__13174),
            .I(N__13168));
    LocalMux I__2258 (
            .O(N__13171),
            .I(N__13165));
    Span4Mux_h I__2257 (
            .O(N__13168),
            .I(N__13162));
    Odrv12 I__2256 (
            .O(N__13165),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    Odrv4 I__2255 (
            .O(N__13162),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    InMux I__2254 (
            .O(N__13157),
            .I(N__13135));
    InMux I__2253 (
            .O(N__13156),
            .I(N__13135));
    InMux I__2252 (
            .O(N__13155),
            .I(N__13135));
    InMux I__2251 (
            .O(N__13154),
            .I(N__13135));
    InMux I__2250 (
            .O(N__13153),
            .I(N__13135));
    InMux I__2249 (
            .O(N__13152),
            .I(N__13135));
    InMux I__2248 (
            .O(N__13151),
            .I(N__13135));
    InMux I__2247 (
            .O(N__13150),
            .I(N__13128));
    LocalMux I__2246 (
            .O(N__13135),
            .I(N__13125));
    InMux I__2245 (
            .O(N__13134),
            .I(N__13120));
    InMux I__2244 (
            .O(N__13133),
            .I(N__13120));
    InMux I__2243 (
            .O(N__13132),
            .I(N__13115));
    InMux I__2242 (
            .O(N__13131),
            .I(N__13115));
    LocalMux I__2241 (
            .O(N__13128),
            .I(N__13110));
    Span4Mux_h I__2240 (
            .O(N__13125),
            .I(N__13110));
    LocalMux I__2239 (
            .O(N__13120),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__2238 (
            .O(N__13115),
            .I(\Lab_UT.di_Stens_1 ));
    Odrv4 I__2237 (
            .O(N__13110),
            .I(\Lab_UT.di_Stens_1 ));
    CascadeMux I__2236 (
            .O(N__13103),
            .I(N__13097));
    CascadeMux I__2235 (
            .O(N__13102),
            .I(N__13094));
    CascadeMux I__2234 (
            .O(N__13101),
            .I(N__13090));
    CascadeMux I__2233 (
            .O(N__13100),
            .I(N__13086));
    InMux I__2232 (
            .O(N__13097),
            .I(N__13069));
    InMux I__2231 (
            .O(N__13094),
            .I(N__13069));
    InMux I__2230 (
            .O(N__13093),
            .I(N__13069));
    InMux I__2229 (
            .O(N__13090),
            .I(N__13069));
    InMux I__2228 (
            .O(N__13089),
            .I(N__13069));
    InMux I__2227 (
            .O(N__13086),
            .I(N__13069));
    InMux I__2226 (
            .O(N__13085),
            .I(N__13069));
    InMux I__2225 (
            .O(N__13084),
            .I(N__13065));
    LocalMux I__2224 (
            .O(N__13069),
            .I(N__13058));
    InMux I__2223 (
            .O(N__13068),
            .I(N__13055));
    LocalMux I__2222 (
            .O(N__13065),
            .I(N__13052));
    InMux I__2221 (
            .O(N__13064),
            .I(N__13049));
    InMux I__2220 (
            .O(N__13063),
            .I(N__13046));
    InMux I__2219 (
            .O(N__13062),
            .I(N__13041));
    InMux I__2218 (
            .O(N__13061),
            .I(N__13041));
    Span4Mux_h I__2217 (
            .O(N__13058),
            .I(N__13038));
    LocalMux I__2216 (
            .O(N__13055),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv12 I__2215 (
            .O(N__13052),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2214 (
            .O(N__13049),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2213 (
            .O(N__13046),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2212 (
            .O(N__13041),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv4 I__2211 (
            .O(N__13038),
            .I(\Lab_UT.di_Stens_0 ));
    CascadeMux I__2210 (
            .O(N__13025),
            .I(N__13019));
    CascadeMux I__2209 (
            .O(N__13024),
            .I(N__13014));
    CascadeMux I__2208 (
            .O(N__13023),
            .I(N__13010));
    CascadeMux I__2207 (
            .O(N__13022),
            .I(N__13006));
    InMux I__2206 (
            .O(N__13019),
            .I(N__13001));
    InMux I__2205 (
            .O(N__13018),
            .I(N__12986));
    InMux I__2204 (
            .O(N__13017),
            .I(N__12986));
    InMux I__2203 (
            .O(N__13014),
            .I(N__12986));
    InMux I__2202 (
            .O(N__13013),
            .I(N__12986));
    InMux I__2201 (
            .O(N__13010),
            .I(N__12986));
    InMux I__2200 (
            .O(N__13009),
            .I(N__12986));
    InMux I__2199 (
            .O(N__13006),
            .I(N__12986));
    InMux I__2198 (
            .O(N__13005),
            .I(N__12981));
    InMux I__2197 (
            .O(N__13004),
            .I(N__12981));
    LocalMux I__2196 (
            .O(N__13001),
            .I(N__12976));
    LocalMux I__2195 (
            .O(N__12986),
            .I(N__12976));
    LocalMux I__2194 (
            .O(N__12981),
            .I(\Lab_UT.di_Stens_3 ));
    Odrv4 I__2193 (
            .O(N__12976),
            .I(\Lab_UT.di_Stens_3 ));
    InMux I__2192 (
            .O(N__12971),
            .I(N__12960));
    InMux I__2191 (
            .O(N__12970),
            .I(N__12954));
    InMux I__2190 (
            .O(N__12969),
            .I(N__12939));
    InMux I__2189 (
            .O(N__12968),
            .I(N__12939));
    InMux I__2188 (
            .O(N__12967),
            .I(N__12939));
    InMux I__2187 (
            .O(N__12966),
            .I(N__12939));
    InMux I__2186 (
            .O(N__12965),
            .I(N__12939));
    InMux I__2185 (
            .O(N__12964),
            .I(N__12939));
    InMux I__2184 (
            .O(N__12963),
            .I(N__12939));
    LocalMux I__2183 (
            .O(N__12960),
            .I(N__12936));
    InMux I__2182 (
            .O(N__12959),
            .I(N__12933));
    InMux I__2181 (
            .O(N__12958),
            .I(N__12928));
    InMux I__2180 (
            .O(N__12957),
            .I(N__12928));
    LocalMux I__2179 (
            .O(N__12954),
            .I(N__12923));
    LocalMux I__2178 (
            .O(N__12939),
            .I(N__12923));
    Span4Mux_h I__2177 (
            .O(N__12936),
            .I(N__12920));
    LocalMux I__2176 (
            .O(N__12933),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__2175 (
            .O(N__12928),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv4 I__2174 (
            .O(N__12923),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv4 I__2173 (
            .O(N__12920),
            .I(\Lab_UT.di_Stens_2 ));
    InMux I__2172 (
            .O(N__12911),
            .I(N__12908));
    LocalMux I__2171 (
            .O(N__12908),
            .I(\Lab_UT.didp.countrce3.q_5_3 ));
    CascadeMux I__2170 (
            .O(N__12905),
            .I(N__12901));
    CascadeMux I__2169 (
            .O(N__12904),
            .I(N__12898));
    InMux I__2168 (
            .O(N__12901),
            .I(N__12895));
    InMux I__2167 (
            .O(N__12898),
            .I(N__12892));
    LocalMux I__2166 (
            .O(N__12895),
            .I(\Lab_UT.didp.q_fast_1 ));
    LocalMux I__2165 (
            .O(N__12892),
            .I(\Lab_UT.didp.q_fast_1 ));
    InMux I__2164 (
            .O(N__12887),
            .I(N__12884));
    LocalMux I__2163 (
            .O(N__12884),
            .I(\Lab_UT.didp.countrce4.q_5_1 ));
    CascadeMux I__2162 (
            .O(N__12881),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__2161 (
            .O(N__12878),
            .I(N__12875));
    LocalMux I__2160 (
            .O(N__12875),
            .I(N__12871));
    CascadeMux I__2159 (
            .O(N__12874),
            .I(N__12868));
    Span4Mux_h I__2158 (
            .O(N__12871),
            .I(N__12864));
    InMux I__2157 (
            .O(N__12868),
            .I(N__12859));
    InMux I__2156 (
            .O(N__12867),
            .I(N__12859));
    Odrv4 I__2155 (
            .O(N__12864),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_0 ));
    LocalMux I__2154 (
            .O(N__12859),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_0 ));
    InMux I__2153 (
            .O(N__12854),
            .I(N__12845));
    InMux I__2152 (
            .O(N__12853),
            .I(N__12845));
    InMux I__2151 (
            .O(N__12852),
            .I(N__12840));
    InMux I__2150 (
            .O(N__12851),
            .I(N__12840));
    InMux I__2149 (
            .O(N__12850),
            .I(N__12837));
    LocalMux I__2148 (
            .O(N__12845),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    LocalMux I__2147 (
            .O(N__12840),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    LocalMux I__2146 (
            .O(N__12837),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    CascadeMux I__2145 (
            .O(N__12830),
            .I(N__12824));
    InMux I__2144 (
            .O(N__12829),
            .I(N__12816));
    InMux I__2143 (
            .O(N__12828),
            .I(N__12816));
    InMux I__2142 (
            .O(N__12827),
            .I(N__12816));
    InMux I__2141 (
            .O(N__12824),
            .I(N__12811));
    InMux I__2140 (
            .O(N__12823),
            .I(N__12811));
    LocalMux I__2139 (
            .O(N__12816),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ));
    LocalMux I__2138 (
            .O(N__12811),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ));
    InMux I__2137 (
            .O(N__12806),
            .I(N__12795));
    InMux I__2136 (
            .O(N__12805),
            .I(N__12795));
    InMux I__2135 (
            .O(N__12804),
            .I(N__12795));
    InMux I__2134 (
            .O(N__12803),
            .I(N__12790));
    InMux I__2133 (
            .O(N__12802),
            .I(N__12790));
    LocalMux I__2132 (
            .O(N__12795),
            .I(\Lab_UT.dictrl.next_alarmstate_1_1 ));
    LocalMux I__2131 (
            .O(N__12790),
            .I(\Lab_UT.dictrl.next_alarmstate_1_1 ));
    InMux I__2130 (
            .O(N__12785),
            .I(N__12782));
    LocalMux I__2129 (
            .O(N__12782),
            .I(N__12778));
    CascadeMux I__2128 (
            .O(N__12781),
            .I(N__12774));
    Span4Mux_h I__2127 (
            .O(N__12778),
            .I(N__12770));
    InMux I__2126 (
            .O(N__12777),
            .I(N__12767));
    InMux I__2125 (
            .O(N__12774),
            .I(N__12762));
    InMux I__2124 (
            .O(N__12773),
            .I(N__12762));
    Odrv4 I__2123 (
            .O(N__12770),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__2122 (
            .O(N__12767),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__2121 (
            .O(N__12762),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    InMux I__2120 (
            .O(N__12755),
            .I(N__12749));
    InMux I__2119 (
            .O(N__12754),
            .I(N__12749));
    LocalMux I__2118 (
            .O(N__12749),
            .I(N__12746));
    Span4Mux_h I__2117 (
            .O(N__12746),
            .I(N__12739));
    InMux I__2116 (
            .O(N__12745),
            .I(N__12736));
    InMux I__2115 (
            .O(N__12744),
            .I(N__12729));
    InMux I__2114 (
            .O(N__12743),
            .I(N__12729));
    InMux I__2113 (
            .O(N__12742),
            .I(N__12729));
    Odrv4 I__2112 (
            .O(N__12739),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    LocalMux I__2111 (
            .O(N__12736),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    LocalMux I__2110 (
            .O(N__12729),
            .I(\Lab_UT.dictrl.alarmstateZ0Z_1 ));
    InMux I__2109 (
            .O(N__12722),
            .I(N__12719));
    LocalMux I__2108 (
            .O(N__12719),
            .I(\Lab_UT.alarmchar_2_1_1 ));
    InMux I__2107 (
            .O(N__12716),
            .I(N__12713));
    LocalMux I__2106 (
            .O(N__12713),
            .I(N__12708));
    InMux I__2105 (
            .O(N__12712),
            .I(N__12705));
    InMux I__2104 (
            .O(N__12711),
            .I(N__12702));
    Odrv4 I__2103 (
            .O(N__12708),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__2102 (
            .O(N__12705),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__2101 (
            .O(N__12702),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__2100 (
            .O(N__12695),
            .I(N__12689));
    InMux I__2099 (
            .O(N__12694),
            .I(N__12689));
    LocalMux I__2098 (
            .O(N__12689),
            .I(\Lab_UT.didp.countrce2.q_5_1 ));
    CascadeMux I__2097 (
            .O(N__12686),
            .I(N__12683));
    InMux I__2096 (
            .O(N__12683),
            .I(N__12680));
    LocalMux I__2095 (
            .O(N__12680),
            .I(\Lab_UT.didp.countrce2.q_5_2 ));
    InMux I__2094 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__2093 (
            .O(N__12674),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    IoInMux I__2092 (
            .O(N__12671),
            .I(N__12668));
    LocalMux I__2091 (
            .O(N__12668),
            .I(N__12665));
    IoSpan4Mux I__2090 (
            .O(N__12665),
            .I(N__12661));
    SRMux I__2089 (
            .O(N__12664),
            .I(N__12658));
    Span4Mux_s0_v I__2088 (
            .O(N__12661),
            .I(N__12652));
    LocalMux I__2087 (
            .O(N__12658),
            .I(N__12652));
    InMux I__2086 (
            .O(N__12657),
            .I(N__12649));
    Span4Mux_v I__2085 (
            .O(N__12652),
            .I(N__12645));
    LocalMux I__2084 (
            .O(N__12649),
            .I(N__12642));
    CascadeMux I__2083 (
            .O(N__12648),
            .I(N__12639));
    Span4Mux_v I__2082 (
            .O(N__12645),
            .I(N__12636));
    Span4Mux_v I__2081 (
            .O(N__12642),
            .I(N__12633));
    InMux I__2080 (
            .O(N__12639),
            .I(N__12630));
    Odrv4 I__2079 (
            .O(N__12636),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2078 (
            .O(N__12633),
            .I(CONSTANT_ONE_NET));
    LocalMux I__2077 (
            .O(N__12630),
            .I(CONSTANT_ONE_NET));
    CEMux I__2076 (
            .O(N__12623),
            .I(N__12620));
    LocalMux I__2075 (
            .O(N__12620),
            .I(N__12617));
    Odrv4 I__2074 (
            .O(N__12617),
            .I(\Lab_UT.dictrl.G_64 ));
    InMux I__2073 (
            .O(N__12614),
            .I(N__12608));
    InMux I__2072 (
            .O(N__12613),
            .I(N__12608));
    LocalMux I__2071 (
            .O(N__12608),
            .I(\Lab_UT.alarmMatch ));
    CascadeMux I__2070 (
            .O(N__12605),
            .I(\Lab_UT.dictrl.idle_cascade_ ));
    CascadeMux I__2069 (
            .O(N__12602),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ));
    InMux I__2068 (
            .O(N__12599),
            .I(N__12596));
    LocalMux I__2067 (
            .O(N__12596),
            .I(\Lab_UT.alarmchar9 ));
    InMux I__2066 (
            .O(N__12593),
            .I(N__12590));
    LocalMux I__2065 (
            .O(N__12590),
            .I(N__12587));
    Odrv4 I__2064 (
            .O(N__12587),
            .I(\Lab_UT.alarmchar10 ));
    InMux I__2063 (
            .O(N__12584),
            .I(N__12581));
    LocalMux I__2062 (
            .O(N__12581),
            .I(N__12578));
    Span4Mux_h I__2061 (
            .O(N__12578),
            .I(N__12575));
    Odrv4 I__2060 (
            .O(N__12575),
            .I(\Lab_UT.alarmchar10_i_2 ));
    CascadeMux I__2059 (
            .O(N__12572),
            .I(\Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_ ));
    CascadeMux I__2058 (
            .O(N__12569),
            .I(\uu2.N_57_cascade_ ));
    CascadeMux I__2057 (
            .O(N__12566),
            .I(N__12563));
    InMux I__2056 (
            .O(N__12563),
            .I(N__12557));
    InMux I__2055 (
            .O(N__12562),
            .I(N__12557));
    LocalMux I__2054 (
            .O(N__12557),
            .I(N__12553));
    InMux I__2053 (
            .O(N__12556),
            .I(N__12550));
    Odrv4 I__2052 (
            .O(N__12553),
            .I(\uu2.w_data_i_a3_0_5 ));
    LocalMux I__2051 (
            .O(N__12550),
            .I(\uu2.w_data_i_a3_0_5 ));
    CascadeMux I__2050 (
            .O(N__12545),
            .I(\uu2.mem0.w_data_0_a3_0_6_cascade_ ));
    InMux I__2049 (
            .O(N__12542),
            .I(N__12539));
    LocalMux I__2048 (
            .O(N__12539),
            .I(N__12536));
    Span4Mux_v I__2047 (
            .O(N__12536),
            .I(N__12533));
    Span4Mux_s3_h I__2046 (
            .O(N__12533),
            .I(N__12530));
    Odrv4 I__2045 (
            .O(N__12530),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__2044 (
            .O(N__12527),
            .I(N__12522));
    InMux I__2043 (
            .O(N__12526),
            .I(N__12517));
    InMux I__2042 (
            .O(N__12525),
            .I(N__12517));
    LocalMux I__2041 (
            .O(N__12522),
            .I(\uu2.w_data_displaying_2_i_a2_i_a2_0_0 ));
    LocalMux I__2040 (
            .O(N__12517),
            .I(\uu2.w_data_displaying_2_i_a2_i_a2_0_0 ));
    InMux I__2039 (
            .O(N__12512),
            .I(N__12509));
    LocalMux I__2038 (
            .O(N__12509),
            .I(N__12506));
    Odrv12 I__2037 (
            .O(N__12506),
            .I(\Lab_UT.alarmcharZ0Z_4 ));
    CascadeMux I__2036 (
            .O(N__12503),
            .I(N__12498));
    InMux I__2035 (
            .O(N__12502),
            .I(N__12495));
    InMux I__2034 (
            .O(N__12501),
            .I(N__12492));
    InMux I__2033 (
            .O(N__12498),
            .I(N__12489));
    LocalMux I__2032 (
            .O(N__12495),
            .I(L3_tx_data_6));
    LocalMux I__2031 (
            .O(N__12492),
            .I(L3_tx_data_6));
    LocalMux I__2030 (
            .O(N__12489),
            .I(L3_tx_data_6));
    InMux I__2029 (
            .O(N__12482),
            .I(N__12477));
    InMux I__2028 (
            .O(N__12481),
            .I(N__12472));
    InMux I__2027 (
            .O(N__12480),
            .I(N__12472));
    LocalMux I__2026 (
            .O(N__12477),
            .I(L3_tx_data_3));
    LocalMux I__2025 (
            .O(N__12472),
            .I(L3_tx_data_3));
    InMux I__2024 (
            .O(N__12467),
            .I(N__12464));
    LocalMux I__2023 (
            .O(N__12464),
            .I(N__12459));
    InMux I__2022 (
            .O(N__12463),
            .I(N__12456));
    InMux I__2021 (
            .O(N__12462),
            .I(N__12453));
    Odrv4 I__2020 (
            .O(N__12459),
            .I(L3_tx_data_0));
    LocalMux I__2019 (
            .O(N__12456),
            .I(L3_tx_data_0));
    LocalMux I__2018 (
            .O(N__12453),
            .I(L3_tx_data_0));
    InMux I__2017 (
            .O(N__12446),
            .I(N__12443));
    LocalMux I__2016 (
            .O(N__12443),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    CascadeMux I__2015 (
            .O(N__12440),
            .I(uu2_un1_w_user_cr_0_cascade_));
    CascadeMux I__2014 (
            .O(N__12437),
            .I(N__12433));
    CascadeMux I__2013 (
            .O(N__12436),
            .I(N__12429));
    InMux I__2012 (
            .O(N__12433),
            .I(N__12426));
    InMux I__2011 (
            .O(N__12432),
            .I(N__12421));
    InMux I__2010 (
            .O(N__12429),
            .I(N__12421));
    LocalMux I__2009 (
            .O(N__12426),
            .I(L3_tx_data_2));
    LocalMux I__2008 (
            .O(N__12421),
            .I(L3_tx_data_2));
    InMux I__2007 (
            .O(N__12416),
            .I(N__12413));
    LocalMux I__2006 (
            .O(N__12413),
            .I(N__12410));
    Span4Mux_v I__2005 (
            .O(N__12410),
            .I(N__12407));
    Odrv4 I__2004 (
            .O(N__12407),
            .I(\uu2.mem0.w_data_2 ));
    InMux I__2003 (
            .O(N__12404),
            .I(N__12401));
    LocalMux I__2002 (
            .O(N__12401),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_44 ));
    CascadeMux I__2001 (
            .O(N__12398),
            .I(N__12395));
    InMux I__2000 (
            .O(N__12395),
            .I(N__12392));
    LocalMux I__1999 (
            .O(N__12392),
            .I(N__12389));
    Odrv4 I__1998 (
            .O(N__12389),
            .I(\uu2.mem0.w_addr_2 ));
    CascadeMux I__1997 (
            .O(N__12386),
            .I(\uu2.mem0.bitmap_pmux_sn_N_33_cascade_ ));
    InMux I__1996 (
            .O(N__12383),
            .I(N__12380));
    LocalMux I__1995 (
            .O(N__12380),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ));
    CascadeMux I__1994 (
            .O(N__12377),
            .I(N__12373));
    CascadeMux I__1993 (
            .O(N__12376),
            .I(N__12370));
    InMux I__1992 (
            .O(N__12373),
            .I(N__12367));
    InMux I__1991 (
            .O(N__12370),
            .I(N__12364));
    LocalMux I__1990 (
            .O(N__12367),
            .I(\uu2.N_34 ));
    LocalMux I__1989 (
            .O(N__12364),
            .I(\uu2.N_34 ));
    InMux I__1988 (
            .O(N__12359),
            .I(N__12356));
    LocalMux I__1987 (
            .O(N__12356),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_42 ));
    InMux I__1986 (
            .O(N__12353),
            .I(N__12347));
    InMux I__1985 (
            .O(N__12352),
            .I(N__12347));
    LocalMux I__1984 (
            .O(N__12347),
            .I(N__12344));
    Odrv4 I__1983 (
            .O(N__12344),
            .I(\uu2.N_49 ));
    CascadeMux I__1982 (
            .O(N__12341),
            .I(N__12337));
    InMux I__1981 (
            .O(N__12340),
            .I(N__12334));
    InMux I__1980 (
            .O(N__12337),
            .I(N__12331));
    LocalMux I__1979 (
            .O(N__12334),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__1978 (
            .O(N__12331),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1977 (
            .O(N__12326),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__1976 (
            .O(N__12323),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__1975 (
            .O(N__12320),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__1974 (
            .O(N__12317),
            .I(N__12308));
    InMux I__1973 (
            .O(N__12316),
            .I(N__12308));
    InMux I__1972 (
            .O(N__12315),
            .I(N__12308));
    LocalMux I__1971 (
            .O(N__12308),
            .I(\buart.Z_tx.ser_clk ));
    InMux I__1970 (
            .O(N__12305),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    InMux I__1969 (
            .O(N__12302),
            .I(N__12299));
    LocalMux I__1968 (
            .O(N__12299),
            .I(\uu2.un3_w_addr_user_4 ));
    InMux I__1967 (
            .O(N__12296),
            .I(N__12290));
    InMux I__1966 (
            .O(N__12295),
            .I(N__12290));
    LocalMux I__1965 (
            .O(N__12290),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    InMux I__1964 (
            .O(N__12287),
            .I(N__12281));
    InMux I__1963 (
            .O(N__12286),
            .I(N__12281));
    LocalMux I__1962 (
            .O(N__12281),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1961 (
            .O(N__12278),
            .I(N__12274));
    InMux I__1960 (
            .O(N__12277),
            .I(N__12269));
    InMux I__1959 (
            .O(N__12274),
            .I(N__12269));
    LocalMux I__1958 (
            .O(N__12269),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__1957 (
            .O(N__12266),
            .I(N__12260));
    InMux I__1956 (
            .O(N__12265),
            .I(N__12260));
    LocalMux I__1955 (
            .O(N__12260),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1954 (
            .O(N__12257),
            .I(N__12254));
    LocalMux I__1953 (
            .O(N__12254),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__1952 (
            .O(N__12251),
            .I(N__12248));
    InMux I__1951 (
            .O(N__12248),
            .I(N__12245));
    LocalMux I__1950 (
            .O(N__12245),
            .I(N__12242));
    Span4Mux_s3_h I__1949 (
            .O(N__12242),
            .I(N__12239));
    Odrv4 I__1948 (
            .O(N__12239),
            .I(\uu2.mem0.w_addr_8 ));
    CascadeMux I__1947 (
            .O(N__12236),
            .I(N__12233));
    InMux I__1946 (
            .O(N__12233),
            .I(N__12230));
    LocalMux I__1945 (
            .O(N__12230),
            .I(N__12227));
    Odrv12 I__1944 (
            .O(N__12227),
            .I(\uu2.mem0.w_addr_0 ));
    CascadeMux I__1943 (
            .O(N__12224),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    InMux I__1942 (
            .O(N__12221),
            .I(N__12218));
    LocalMux I__1941 (
            .O(N__12218),
            .I(\buart.Z_rx.un1_sample_0 ));
    CascadeMux I__1940 (
            .O(N__12215),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    InMux I__1939 (
            .O(N__12212),
            .I(N__12209));
    LocalMux I__1938 (
            .O(N__12209),
            .I(N__12202));
    InMux I__1937 (
            .O(N__12208),
            .I(N__12199));
    InMux I__1936 (
            .O(N__12207),
            .I(N__12194));
    InMux I__1935 (
            .O(N__12206),
            .I(N__12194));
    InMux I__1934 (
            .O(N__12205),
            .I(N__12191));
    Span4Mux_v I__1933 (
            .O(N__12202),
            .I(N__12188));
    LocalMux I__1932 (
            .O(N__12199),
            .I(N__12183));
    LocalMux I__1931 (
            .O(N__12194),
            .I(N__12183));
    LocalMux I__1930 (
            .O(N__12191),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv4 I__1929 (
            .O(N__12188),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv12 I__1928 (
            .O(N__12183),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    IoInMux I__1927 (
            .O(N__12176),
            .I(N__12173));
    LocalMux I__1926 (
            .O(N__12173),
            .I(N__12170));
    Span4Mux_s3_v I__1925 (
            .O(N__12170),
            .I(N__12167));
    Odrv4 I__1924 (
            .O(N__12167),
            .I(\buart.Z_rx.sample ));
    InMux I__1923 (
            .O(N__12164),
            .I(N__12160));
    InMux I__1922 (
            .O(N__12163),
            .I(N__12157));
    LocalMux I__1921 (
            .O(N__12160),
            .I(N__12154));
    LocalMux I__1920 (
            .O(N__12157),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv12 I__1919 (
            .O(N__12154),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1918 (
            .O(N__12149),
            .I(N__12143));
    InMux I__1917 (
            .O(N__12148),
            .I(N__12143));
    LocalMux I__1916 (
            .O(N__12143),
            .I(\buart.Z_rx.idle ));
    CascadeMux I__1915 (
            .O(N__12140),
            .I(\buart.Z_rx.startbit_cascade_ ));
    InMux I__1914 (
            .O(N__12137),
            .I(N__12132));
    InMux I__1913 (
            .O(N__12136),
            .I(N__12129));
    InMux I__1912 (
            .O(N__12135),
            .I(N__12126));
    LocalMux I__1911 (
            .O(N__12132),
            .I(bu_rx_data_rdy));
    LocalMux I__1910 (
            .O(N__12129),
            .I(bu_rx_data_rdy));
    LocalMux I__1909 (
            .O(N__12126),
            .I(bu_rx_data_rdy));
    CEMux I__1908 (
            .O(N__12119),
            .I(N__12116));
    LocalMux I__1907 (
            .O(N__12116),
            .I(N__12111));
    CEMux I__1906 (
            .O(N__12115),
            .I(N__12108));
    CEMux I__1905 (
            .O(N__12114),
            .I(N__12105));
    Span4Mux_v I__1904 (
            .O(N__12111),
            .I(N__12100));
    LocalMux I__1903 (
            .O(N__12108),
            .I(N__12100));
    LocalMux I__1902 (
            .O(N__12105),
            .I(N__12097));
    Odrv4 I__1901 (
            .O(N__12100),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__1900 (
            .O(N__12097),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__1899 (
            .O(N__12092),
            .I(N__12086));
    InMux I__1898 (
            .O(N__12091),
            .I(N__12086));
    LocalMux I__1897 (
            .O(N__12086),
            .I(N__12083));
    Span4Mux_v I__1896 (
            .O(N__12083),
            .I(N__12080));
    Odrv4 I__1895 (
            .O(N__12080),
            .I(\Lab_UT.didp.countrce2.q_5_0 ));
    InMux I__1894 (
            .O(N__12077),
            .I(N__12071));
    InMux I__1893 (
            .O(N__12076),
            .I(N__12064));
    InMux I__1892 (
            .O(N__12075),
            .I(N__12064));
    InMux I__1891 (
            .O(N__12074),
            .I(N__12064));
    LocalMux I__1890 (
            .O(N__12071),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1889 (
            .O(N__12064),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1888 (
            .O(N__12059),
            .I(N__12056));
    InMux I__1887 (
            .O(N__12056),
            .I(N__12051));
    InMux I__1886 (
            .O(N__12055),
            .I(N__12046));
    InMux I__1885 (
            .O(N__12054),
            .I(N__12046));
    LocalMux I__1884 (
            .O(N__12051),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1883 (
            .O(N__12046),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1882 (
            .O(N__12041),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    CascadeMux I__1881 (
            .O(N__12038),
            .I(\Lab_UT.dicLdAMones_0_cascade_ ));
    InMux I__1880 (
            .O(N__12035),
            .I(N__12032));
    LocalMux I__1879 (
            .O(N__12032),
            .I(N__12028));
    InMux I__1878 (
            .O(N__12031),
            .I(N__12024));
    Span4Mux_v I__1877 (
            .O(N__12028),
            .I(N__12021));
    InMux I__1876 (
            .O(N__12027),
            .I(N__12018));
    LocalMux I__1875 (
            .O(N__12024),
            .I(N__12015));
    Odrv4 I__1874 (
            .O(N__12021),
            .I(\Lab_UT.di_AMones_0 ));
    LocalMux I__1873 (
            .O(N__12018),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv12 I__1872 (
            .O(N__12015),
            .I(\Lab_UT.di_AMones_0 ));
    InMux I__1871 (
            .O(N__12008),
            .I(N__12005));
    LocalMux I__1870 (
            .O(N__12005),
            .I(N__12000));
    InMux I__1869 (
            .O(N__12004),
            .I(N__11997));
    InMux I__1868 (
            .O(N__12003),
            .I(N__11994));
    Span4Mux_v I__1867 (
            .O(N__12000),
            .I(N__11989));
    LocalMux I__1866 (
            .O(N__11997),
            .I(N__11989));
    LocalMux I__1865 (
            .O(N__11994),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__1864 (
            .O(N__11989),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__1863 (
            .O(N__11984),
            .I(N__11981));
    LocalMux I__1862 (
            .O(N__11981),
            .I(N__11976));
    InMux I__1861 (
            .O(N__11980),
            .I(N__11973));
    InMux I__1860 (
            .O(N__11979),
            .I(N__11970));
    Span4Mux_v I__1859 (
            .O(N__11976),
            .I(N__11965));
    LocalMux I__1858 (
            .O(N__11973),
            .I(N__11965));
    LocalMux I__1857 (
            .O(N__11970),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__1856 (
            .O(N__11965),
            .I(\Lab_UT.di_AMones_2 ));
    CascadeMux I__1855 (
            .O(N__11960),
            .I(N__11956));
    InMux I__1854 (
            .O(N__11959),
            .I(N__11948));
    InMux I__1853 (
            .O(N__11956),
            .I(N__11948));
    InMux I__1852 (
            .O(N__11955),
            .I(N__11948));
    LocalMux I__1851 (
            .O(N__11948),
            .I(\Lab_UT.dicLdAMones_0 ));
    CascadeMux I__1850 (
            .O(N__11945),
            .I(N__11940));
    InMux I__1849 (
            .O(N__11944),
            .I(N__11937));
    InMux I__1848 (
            .O(N__11943),
            .I(N__11934));
    InMux I__1847 (
            .O(N__11940),
            .I(N__11931));
    LocalMux I__1846 (
            .O(N__11937),
            .I(N__11926));
    LocalMux I__1845 (
            .O(N__11934),
            .I(N__11926));
    LocalMux I__1844 (
            .O(N__11931),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__1843 (
            .O(N__11926),
            .I(\Lab_UT.di_AMones_3 ));
    InMux I__1842 (
            .O(N__11921),
            .I(N__11918));
    LocalMux I__1841 (
            .O(N__11918),
            .I(N__11915));
    Span4Mux_v I__1840 (
            .O(N__11915),
            .I(N__11912));
    Odrv4 I__1839 (
            .O(N__11912),
            .I(\resetGen.escKeyZ0Z_5 ));
    CascadeMux I__1838 (
            .O(N__11909),
            .I(\resetGen.escKeyZ0Z_4_cascade_ ));
    CascadeMux I__1837 (
            .O(N__11906),
            .I(\Lab_UT.didp.countrce3.q_5_3_cascade_ ));
    InMux I__1836 (
            .O(N__11903),
            .I(N__11897));
    InMux I__1835 (
            .O(N__11902),
            .I(N__11897));
    LocalMux I__1834 (
            .O(N__11897),
            .I(\Lab_UT.didp.countrce3.q_fastZ0Z_3 ));
    CascadeMux I__1833 (
            .O(N__11894),
            .I(N__11890));
    InMux I__1832 (
            .O(N__11893),
            .I(N__11885));
    InMux I__1831 (
            .O(N__11890),
            .I(N__11885));
    LocalMux I__1830 (
            .O(N__11885),
            .I(\Lab_UT.didp.q_fast_3 ));
    InMux I__1829 (
            .O(N__11882),
            .I(N__11879));
    LocalMux I__1828 (
            .O(N__11879),
            .I(\Lab_UT.didp.countrce3.did_alarmMatch_0 ));
    InMux I__1827 (
            .O(N__11876),
            .I(N__11872));
    InMux I__1826 (
            .O(N__11875),
            .I(N__11869));
    LocalMux I__1825 (
            .O(N__11872),
            .I(N__11866));
    LocalMux I__1824 (
            .O(N__11869),
            .I(N__11863));
    Odrv12 I__1823 (
            .O(N__11866),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__1822 (
            .O(N__11863),
            .I(\Lab_UT.di_AMtens_0 ));
    InMux I__1821 (
            .O(N__11858),
            .I(N__11854));
    InMux I__1820 (
            .O(N__11857),
            .I(N__11851));
    LocalMux I__1819 (
            .O(N__11854),
            .I(N__11848));
    LocalMux I__1818 (
            .O(N__11851),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv4 I__1817 (
            .O(N__11848),
            .I(\Lab_UT.di_AMtens_1 ));
    InMux I__1816 (
            .O(N__11843),
            .I(N__11837));
    InMux I__1815 (
            .O(N__11842),
            .I(N__11837));
    LocalMux I__1814 (
            .O(N__11837),
            .I(N__11834));
    Odrv12 I__1813 (
            .O(N__11834),
            .I(\Lab_UT.di_AMtens_2 ));
    InMux I__1812 (
            .O(N__11831),
            .I(N__11828));
    LocalMux I__1811 (
            .O(N__11828),
            .I(N__11824));
    InMux I__1810 (
            .O(N__11827),
            .I(N__11821));
    Odrv12 I__1809 (
            .O(N__11824),
            .I(\Lab_UT.di_AMtens_3 ));
    LocalMux I__1808 (
            .O(N__11821),
            .I(\Lab_UT.di_AMtens_3 ));
    CascadeMux I__1807 (
            .O(N__11816),
            .I(\Lab_UT.three_2_0_cascade_ ));
    InMux I__1806 (
            .O(N__11813),
            .I(N__11809));
    InMux I__1805 (
            .O(N__11812),
            .I(N__11806));
    LocalMux I__1804 (
            .O(N__11809),
            .I(N__11803));
    LocalMux I__1803 (
            .O(N__11806),
            .I(N__11800));
    Odrv12 I__1802 (
            .O(N__11803),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__1801 (
            .O(N__11800),
            .I(\Lab_UT.di_ASones_1 ));
    InMux I__1800 (
            .O(N__11795),
            .I(N__11792));
    LocalMux I__1799 (
            .O(N__11792),
            .I(\Lab_UT.didp.did_alarmMatch_3 ));
    CascadeMux I__1798 (
            .O(N__11789),
            .I(N__11786));
    InMux I__1797 (
            .O(N__11786),
            .I(N__11782));
    InMux I__1796 (
            .O(N__11785),
            .I(N__11779));
    LocalMux I__1795 (
            .O(N__11782),
            .I(\Lab_UT.didp.countrce2.q_fastZ0Z_1 ));
    LocalMux I__1794 (
            .O(N__11779),
            .I(\Lab_UT.didp.countrce2.q_fastZ0Z_1 ));
    InMux I__1793 (
            .O(N__11774),
            .I(N__11770));
    InMux I__1792 (
            .O(N__11773),
            .I(N__11767));
    LocalMux I__1791 (
            .O(N__11770),
            .I(\Lab_UT.didp.countrce3.q_fastZ0Z_1 ));
    LocalMux I__1790 (
            .O(N__11767),
            .I(\Lab_UT.didp.countrce3.q_fastZ0Z_1 ));
    CascadeMux I__1789 (
            .O(N__11762),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    CascadeMux I__1788 (
            .O(N__11759),
            .I(N__11756));
    InMux I__1787 (
            .O(N__11756),
            .I(N__11752));
    InMux I__1786 (
            .O(N__11755),
            .I(N__11748));
    LocalMux I__1785 (
            .O(N__11752),
            .I(N__11745));
    InMux I__1784 (
            .O(N__11751),
            .I(N__11742));
    LocalMux I__1783 (
            .O(N__11748),
            .I(N__11739));
    Odrv4 I__1782 (
            .O(N__11745),
            .I(\Lab_UT.didp.q_fast_0 ));
    LocalMux I__1781 (
            .O(N__11742),
            .I(\Lab_UT.didp.q_fast_0 ));
    Odrv4 I__1780 (
            .O(N__11739),
            .I(\Lab_UT.didp.q_fast_0 ));
    InMux I__1779 (
            .O(N__11732),
            .I(N__11729));
    LocalMux I__1778 (
            .O(N__11729),
            .I(N__11726));
    Odrv4 I__1777 (
            .O(N__11726),
            .I(\Lab_UT.didp.countrce2.un20_qPone ));
    CascadeMux I__1776 (
            .O(N__11723),
            .I(\Lab_UT.didp.countrce2.q_5_3_cascade_ ));
    InMux I__1775 (
            .O(N__11720),
            .I(N__11717));
    LocalMux I__1774 (
            .O(N__11717),
            .I(N__11712));
    InMux I__1773 (
            .O(N__11716),
            .I(N__11709));
    InMux I__1772 (
            .O(N__11715),
            .I(N__11706));
    Odrv4 I__1771 (
            .O(N__11712),
            .I(\Lab_UT.di_AStens_3 ));
    LocalMux I__1770 (
            .O(N__11709),
            .I(\Lab_UT.di_AStens_3 ));
    LocalMux I__1769 (
            .O(N__11706),
            .I(\Lab_UT.di_AStens_3 ));
    InMux I__1768 (
            .O(N__11699),
            .I(N__11696));
    LocalMux I__1767 (
            .O(N__11696),
            .I(N__11692));
    InMux I__1766 (
            .O(N__11695),
            .I(N__11689));
    Odrv4 I__1765 (
            .O(N__11692),
            .I(\Lab_UT.didp.countrce2.q_fastZ0Z_3 ));
    LocalMux I__1764 (
            .O(N__11689),
            .I(\Lab_UT.didp.countrce2.q_fastZ0Z_3 ));
    InMux I__1763 (
            .O(N__11684),
            .I(N__11680));
    InMux I__1762 (
            .O(N__11683),
            .I(N__11677));
    LocalMux I__1761 (
            .O(N__11680),
            .I(N__11674));
    LocalMux I__1760 (
            .O(N__11677),
            .I(N__11671));
    Span4Mux_v I__1759 (
            .O(N__11674),
            .I(N__11668));
    Span4Mux_h I__1758 (
            .O(N__11671),
            .I(N__11665));
    Odrv4 I__1757 (
            .O(N__11668),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__1756 (
            .O(N__11665),
            .I(\Lab_UT.di_ASones_3 ));
    InMux I__1755 (
            .O(N__11660),
            .I(N__11657));
    LocalMux I__1754 (
            .O(N__11657),
            .I(\Lab_UT.didp.countrce2.q_5_3 ));
    InMux I__1753 (
            .O(N__11654),
            .I(N__11651));
    LocalMux I__1752 (
            .O(N__11651),
            .I(\Lab_UT.didp.did_alarmMatch_2 ));
    CascadeMux I__1751 (
            .O(N__11648),
            .I(\Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_ ));
    InMux I__1750 (
            .O(N__11645),
            .I(N__11642));
    LocalMux I__1749 (
            .O(N__11642),
            .I(\Lab_UT.didp.did_alarmMatch_12 ));
    InMux I__1748 (
            .O(N__11639),
            .I(N__11636));
    LocalMux I__1747 (
            .O(N__11636),
            .I(\Lab_UT.min1Z0Z_0 ));
    InMux I__1746 (
            .O(N__11633),
            .I(N__11630));
    LocalMux I__1745 (
            .O(N__11630),
            .I(N__11627));
    Odrv4 I__1744 (
            .O(N__11627),
            .I(\Lab_UT.dispString.m25_ns_1 ));
    CascadeMux I__1743 (
            .O(N__11624),
            .I(N__11621));
    InMux I__1742 (
            .O(N__11621),
            .I(N__11618));
    LocalMux I__1741 (
            .O(N__11618),
            .I(\Lab_UT.min1Z0Z_2 ));
    InMux I__1740 (
            .O(N__11615),
            .I(N__11612));
    LocalMux I__1739 (
            .O(N__11612),
            .I(N__11609));
    Odrv12 I__1738 (
            .O(N__11609),
            .I(\Lab_UT.dispString.N_65 ));
    InMux I__1737 (
            .O(N__11606),
            .I(N__11603));
    LocalMux I__1736 (
            .O(N__11603),
            .I(\Lab_UT.alarmcharZ0Z_6 ));
    InMux I__1735 (
            .O(N__11600),
            .I(N__11597));
    LocalMux I__1734 (
            .O(N__11597),
            .I(N__11579));
    InMux I__1733 (
            .O(N__11596),
            .I(N__11574));
    InMux I__1732 (
            .O(N__11595),
            .I(N__11574));
    InMux I__1731 (
            .O(N__11594),
            .I(N__11571));
    InMux I__1730 (
            .O(N__11593),
            .I(N__11564));
    InMux I__1729 (
            .O(N__11592),
            .I(N__11564));
    InMux I__1728 (
            .O(N__11591),
            .I(N__11564));
    InMux I__1727 (
            .O(N__11590),
            .I(N__11555));
    InMux I__1726 (
            .O(N__11589),
            .I(N__11555));
    InMux I__1725 (
            .O(N__11588),
            .I(N__11555));
    InMux I__1724 (
            .O(N__11587),
            .I(N__11555));
    InMux I__1723 (
            .O(N__11586),
            .I(N__11548));
    InMux I__1722 (
            .O(N__11585),
            .I(N__11548));
    InMux I__1721 (
            .O(N__11584),
            .I(N__11548));
    InMux I__1720 (
            .O(N__11583),
            .I(N__11544));
    InMux I__1719 (
            .O(N__11582),
            .I(N__11541));
    Span4Mux_h I__1718 (
            .O(N__11579),
            .I(N__11536));
    LocalMux I__1717 (
            .O(N__11574),
            .I(N__11536));
    LocalMux I__1716 (
            .O(N__11571),
            .I(N__11527));
    LocalMux I__1715 (
            .O(N__11564),
            .I(N__11527));
    LocalMux I__1714 (
            .O(N__11555),
            .I(N__11527));
    LocalMux I__1713 (
            .O(N__11548),
            .I(N__11527));
    InMux I__1712 (
            .O(N__11547),
            .I(N__11524));
    LocalMux I__1711 (
            .O(N__11544),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__1710 (
            .O(N__11541),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__1709 (
            .O(N__11536),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv12 I__1708 (
            .O(N__11527),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__1707 (
            .O(N__11524),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    InMux I__1706 (
            .O(N__11513),
            .I(N__11510));
    LocalMux I__1705 (
            .O(N__11510),
            .I(\Lab_UT.alarmcharZ0Z_2 ));
    CascadeMux I__1704 (
            .O(N__11507),
            .I(N__11504));
    InMux I__1703 (
            .O(N__11504),
            .I(N__11501));
    LocalMux I__1702 (
            .O(N__11501),
            .I(N__11498));
    Span4Mux_h I__1701 (
            .O(N__11498),
            .I(N__11495));
    Odrv4 I__1700 (
            .O(N__11495),
            .I(\Lab_UT.sec2Z0Z_2 ));
    CascadeMux I__1699 (
            .O(N__11492),
            .I(N__11486));
    CascadeMux I__1698 (
            .O(N__11491),
            .I(N__11483));
    InMux I__1697 (
            .O(N__11490),
            .I(N__11465));
    InMux I__1696 (
            .O(N__11489),
            .I(N__11465));
    InMux I__1695 (
            .O(N__11486),
            .I(N__11460));
    InMux I__1694 (
            .O(N__11483),
            .I(N__11460));
    InMux I__1693 (
            .O(N__11482),
            .I(N__11457));
    InMux I__1692 (
            .O(N__11481),
            .I(N__11450));
    InMux I__1691 (
            .O(N__11480),
            .I(N__11450));
    InMux I__1690 (
            .O(N__11479),
            .I(N__11450));
    InMux I__1689 (
            .O(N__11478),
            .I(N__11443));
    InMux I__1688 (
            .O(N__11477),
            .I(N__11443));
    InMux I__1687 (
            .O(N__11476),
            .I(N__11443));
    InMux I__1686 (
            .O(N__11475),
            .I(N__11438));
    InMux I__1685 (
            .O(N__11474),
            .I(N__11431));
    InMux I__1684 (
            .O(N__11473),
            .I(N__11431));
    InMux I__1683 (
            .O(N__11472),
            .I(N__11431));
    InMux I__1682 (
            .O(N__11471),
            .I(N__11426));
    InMux I__1681 (
            .O(N__11470),
            .I(N__11426));
    LocalMux I__1680 (
            .O(N__11465),
            .I(N__11423));
    LocalMux I__1679 (
            .O(N__11460),
            .I(N__11418));
    LocalMux I__1678 (
            .O(N__11457),
            .I(N__11418));
    LocalMux I__1677 (
            .O(N__11450),
            .I(N__11415));
    LocalMux I__1676 (
            .O(N__11443),
            .I(N__11412));
    InMux I__1675 (
            .O(N__11442),
            .I(N__11407));
    InMux I__1674 (
            .O(N__11441),
            .I(N__11407));
    LocalMux I__1673 (
            .O(N__11438),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__1672 (
            .O(N__11431),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__1671 (
            .O(N__11426),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__1670 (
            .O(N__11423),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__1669 (
            .O(N__11418),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__1668 (
            .O(N__11415),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__1667 (
            .O(N__11412),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__1666 (
            .O(N__11407),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    InMux I__1665 (
            .O(N__11390),
            .I(N__11387));
    LocalMux I__1664 (
            .O(N__11387),
            .I(\Lab_UT.dispString.N_68 ));
    InMux I__1663 (
            .O(N__11384),
            .I(N__11381));
    LocalMux I__1662 (
            .O(N__11381),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_5 ));
    InMux I__1661 (
            .O(N__11378),
            .I(N__11375));
    LocalMux I__1660 (
            .O(N__11375),
            .I(N__11372));
    Odrv4 I__1659 (
            .O(N__11372),
            .I(\Lab_UT.didp.did_alarmMatch_11 ));
    CascadeMux I__1658 (
            .O(N__11369),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ));
    CascadeMux I__1657 (
            .O(N__11366),
            .I(\Lab_UT.dispString.N_86_cascade_ ));
    InMux I__1656 (
            .O(N__11363),
            .I(N__11360));
    LocalMux I__1655 (
            .O(N__11360),
            .I(N__11357));
    Odrv4 I__1654 (
            .O(N__11357),
            .I(\Lab_UT.dispString.N_89 ));
    InMux I__1653 (
            .O(N__11354),
            .I(N__11351));
    LocalMux I__1652 (
            .O(N__11351),
            .I(\Lab_UT.min2Z0Z_0 ));
    InMux I__1651 (
            .O(N__11348),
            .I(N__11345));
    LocalMux I__1650 (
            .O(N__11345),
            .I(\Lab_UT.dispString.m49_ns_1 ));
    CascadeMux I__1649 (
            .O(N__11342),
            .I(N__11339));
    InMux I__1648 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1647 (
            .O(N__11336),
            .I(\Lab_UT.sec1Z0Z_0 ));
    CascadeMux I__1646 (
            .O(N__11333),
            .I(N__11322));
    CascadeMux I__1645 (
            .O(N__11332),
            .I(N__11318));
    InMux I__1644 (
            .O(N__11331),
            .I(N__11315));
    InMux I__1643 (
            .O(N__11330),
            .I(N__11308));
    InMux I__1642 (
            .O(N__11329),
            .I(N__11308));
    InMux I__1641 (
            .O(N__11328),
            .I(N__11308));
    InMux I__1640 (
            .O(N__11327),
            .I(N__11305));
    InMux I__1639 (
            .O(N__11326),
            .I(N__11300));
    InMux I__1638 (
            .O(N__11325),
            .I(N__11300));
    InMux I__1637 (
            .O(N__11322),
            .I(N__11297));
    InMux I__1636 (
            .O(N__11321),
            .I(N__11292));
    InMux I__1635 (
            .O(N__11318),
            .I(N__11292));
    LocalMux I__1634 (
            .O(N__11315),
            .I(N__11287));
    LocalMux I__1633 (
            .O(N__11308),
            .I(N__11287));
    LocalMux I__1632 (
            .O(N__11305),
            .I(N__11282));
    LocalMux I__1631 (
            .O(N__11300),
            .I(N__11282));
    LocalMux I__1630 (
            .O(N__11297),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    LocalMux I__1629 (
            .O(N__11292),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__1628 (
            .O(N__11287),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__1627 (
            .O(N__11282),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    InMux I__1626 (
            .O(N__11273),
            .I(N__11270));
    LocalMux I__1625 (
            .O(N__11270),
            .I(N__11265));
    InMux I__1624 (
            .O(N__11269),
            .I(N__11262));
    InMux I__1623 (
            .O(N__11268),
            .I(N__11259));
    Odrv4 I__1622 (
            .O(N__11265),
            .I(L3_tx_data_5));
    LocalMux I__1621 (
            .O(N__11262),
            .I(L3_tx_data_5));
    LocalMux I__1620 (
            .O(N__11259),
            .I(L3_tx_data_5));
    CascadeMux I__1619 (
            .O(N__11252),
            .I(N__11249));
    InMux I__1618 (
            .O(N__11249),
            .I(N__11246));
    LocalMux I__1617 (
            .O(N__11246),
            .I(N__11241));
    InMux I__1616 (
            .O(N__11245),
            .I(N__11238));
    InMux I__1615 (
            .O(N__11244),
            .I(N__11235));
    Odrv4 I__1614 (
            .O(N__11241),
            .I(L3_tx_data_4));
    LocalMux I__1613 (
            .O(N__11238),
            .I(L3_tx_data_4));
    LocalMux I__1612 (
            .O(N__11235),
            .I(L3_tx_data_4));
    CascadeMux I__1611 (
            .O(N__11228),
            .I(N__11224));
    InMux I__1610 (
            .O(N__11227),
            .I(N__11221));
    InMux I__1609 (
            .O(N__11224),
            .I(N__11218));
    LocalMux I__1608 (
            .O(N__11221),
            .I(N__11215));
    LocalMux I__1607 (
            .O(N__11218),
            .I(N__11212));
    Odrv4 I__1606 (
            .O(N__11215),
            .I(\Lab_UT.alarmcharZ0Z_1 ));
    Odrv4 I__1605 (
            .O(N__11212),
            .I(\Lab_UT.alarmcharZ0Z_1 ));
    CascadeMux I__1604 (
            .O(N__11207),
            .I(N__11204));
    InMux I__1603 (
            .O(N__11204),
            .I(N__11201));
    LocalMux I__1602 (
            .O(N__11201),
            .I(N__11198));
    Span4Mux_v I__1601 (
            .O(N__11198),
            .I(N__11195));
    Odrv4 I__1600 (
            .O(N__11195),
            .I(\uu2.mem0.w_addr_3 ));
    InMux I__1599 (
            .O(N__11192),
            .I(N__11189));
    LocalMux I__1598 (
            .O(N__11189),
            .I(\Lab_UT.dispString.m40_ns_1 ));
    CascadeMux I__1597 (
            .O(N__11186),
            .I(N__11183));
    InMux I__1596 (
            .O(N__11183),
            .I(N__11180));
    LocalMux I__1595 (
            .O(N__11180),
            .I(\Lab_UT.min1Z0Z_3 ));
    CascadeMux I__1594 (
            .O(N__11177),
            .I(\Lab_UT.dispString.N_77_cascade_ ));
    InMux I__1593 (
            .O(N__11174),
            .I(N__11171));
    LocalMux I__1592 (
            .O(N__11171),
            .I(\Lab_UT.dispString.N_80 ));
    InMux I__1591 (
            .O(N__11168),
            .I(N__11165));
    LocalMux I__1590 (
            .O(N__11165),
            .I(\Lab_UT.sec2Z0Z_3 ));
    CascadeMux I__1589 (
            .O(N__11162),
            .I(\uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_ ));
    InMux I__1588 (
            .O(N__11159),
            .I(N__11156));
    LocalMux I__1587 (
            .O(N__11156),
            .I(\uu2.mem0.w_data_0_1_3 ));
    CascadeMux I__1586 (
            .O(N__11153),
            .I(N__11150));
    InMux I__1585 (
            .O(N__11150),
            .I(N__11147));
    LocalMux I__1584 (
            .O(N__11147),
            .I(N__11144));
    Odrv12 I__1583 (
            .O(N__11144),
            .I(\uu2.mem0.w_addr_5 ));
    InMux I__1582 (
            .O(N__11141),
            .I(N__11138));
    LocalMux I__1581 (
            .O(N__11138),
            .I(\uu2.mem0.bitmap_pmux_sn_N_33_0 ));
    CascadeMux I__1580 (
            .O(N__11135),
            .I(\uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_ ));
    CascadeMux I__1579 (
            .O(N__11132),
            .I(\uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_ ));
    InMux I__1578 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__1577 (
            .O(N__11126),
            .I(\uu2.mem0.N_409 ));
    CascadeMux I__1576 (
            .O(N__11123),
            .I(\uu2.N_34_cascade_ ));
    CascadeMux I__1575 (
            .O(N__11120),
            .I(N__11117));
    InMux I__1574 (
            .O(N__11117),
            .I(N__11113));
    InMux I__1573 (
            .O(N__11116),
            .I(N__11110));
    LocalMux I__1572 (
            .O(N__11113),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__1571 (
            .O(N__11110),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__1570 (
            .O(N__11105),
            .I(\buart.Z_tx.ser_clk_cascade_ ));
    InMux I__1569 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__1568 (
            .O(N__11099),
            .I(\buart.Z_tx.uart_busy_0_0 ));
    InMux I__1567 (
            .O(N__11096),
            .I(N__11093));
    LocalMux I__1566 (
            .O(N__11093),
            .I(N__11087));
    InMux I__1565 (
            .O(N__11092),
            .I(N__11084));
    InMux I__1564 (
            .O(N__11091),
            .I(N__11078));
    InMux I__1563 (
            .O(N__11090),
            .I(N__11078));
    Span4Mux_v I__1562 (
            .O(N__11087),
            .I(N__11073));
    LocalMux I__1561 (
            .O(N__11084),
            .I(N__11073));
    InMux I__1560 (
            .O(N__11083),
            .I(N__11070));
    LocalMux I__1559 (
            .O(N__11078),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    Odrv4 I__1558 (
            .O(N__11073),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__1557 (
            .O(N__11070),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    CascadeMux I__1556 (
            .O(N__11063),
            .I(N__11059));
    InMux I__1555 (
            .O(N__11062),
            .I(N__11051));
    InMux I__1554 (
            .O(N__11059),
            .I(N__11051));
    InMux I__1553 (
            .O(N__11058),
            .I(N__11051));
    LocalMux I__1552 (
            .O(N__11051),
            .I(N__11047));
    InMux I__1551 (
            .O(N__11050),
            .I(N__11044));
    Span4Mux_v I__1550 (
            .O(N__11047),
            .I(N__11041));
    LocalMux I__1549 (
            .O(N__11044),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    Odrv4 I__1548 (
            .O(N__11041),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__1547 (
            .O(N__11036),
            .I(N__11032));
    InMux I__1546 (
            .O(N__11035),
            .I(N__11026));
    LocalMux I__1545 (
            .O(N__11032),
            .I(N__11023));
    InMux I__1544 (
            .O(N__11031),
            .I(N__11020));
    InMux I__1543 (
            .O(N__11030),
            .I(N__11015));
    InMux I__1542 (
            .O(N__11029),
            .I(N__11015));
    LocalMux I__1541 (
            .O(N__11026),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    Odrv12 I__1540 (
            .O(N__11023),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1539 (
            .O(N__11020),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1538 (
            .O(N__11015),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__1537 (
            .O(N__11006),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    InMux I__1536 (
            .O(N__11003),
            .I(N__10994));
    InMux I__1535 (
            .O(N__11002),
            .I(N__10994));
    InMux I__1534 (
            .O(N__11001),
            .I(N__10994));
    LocalMux I__1533 (
            .O(N__10994),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    InMux I__1532 (
            .O(N__10991),
            .I(N__10988));
    LocalMux I__1531 (
            .O(N__10988),
            .I(\buart.Z_tx.un1_bitcount_c3 ));
    CascadeMux I__1530 (
            .O(N__10985),
            .I(N__10982));
    InMux I__1529 (
            .O(N__10982),
            .I(N__10979));
    LocalMux I__1528 (
            .O(N__10979),
            .I(N__10976));
    Odrv4 I__1527 (
            .O(N__10976),
            .I(\uu2.mem0.w_addr_1 ));
    IoInMux I__1526 (
            .O(N__10973),
            .I(N__10970));
    LocalMux I__1525 (
            .O(N__10970),
            .I(N__10966));
    InMux I__1524 (
            .O(N__10969),
            .I(N__10963));
    Span12Mux_s9_v I__1523 (
            .O(N__10966),
            .I(N__10960));
    LocalMux I__1522 (
            .O(N__10963),
            .I(N__10957));
    Odrv12 I__1521 (
            .O(N__10960),
            .I(clk));
    Odrv4 I__1520 (
            .O(N__10957),
            .I(clk));
    CEMux I__1519 (
            .O(N__10952),
            .I(N__10949));
    LocalMux I__1518 (
            .O(N__10949),
            .I(N__10945));
    SRMux I__1517 (
            .O(N__10948),
            .I(N__10942));
    Span4Mux_h I__1516 (
            .O(N__10945),
            .I(N__10939));
    LocalMux I__1515 (
            .O(N__10942),
            .I(N__10934));
    Span4Mux_s1_h I__1514 (
            .O(N__10939),
            .I(N__10934));
    Odrv4 I__1513 (
            .O(N__10934),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1512 (
            .O(N__10931),
            .I(N__10928));
    InMux I__1511 (
            .O(N__10928),
            .I(N__10925));
    LocalMux I__1510 (
            .O(N__10925),
            .I(N__10922));
    Odrv4 I__1509 (
            .O(N__10922),
            .I(\uu2.mem0.w_addr_4 ));
    InMux I__1508 (
            .O(N__10919),
            .I(N__10912));
    InMux I__1507 (
            .O(N__10918),
            .I(N__10903));
    InMux I__1506 (
            .O(N__10917),
            .I(N__10903));
    InMux I__1505 (
            .O(N__10916),
            .I(N__10903));
    InMux I__1504 (
            .O(N__10915),
            .I(N__10903));
    LocalMux I__1503 (
            .O(N__10912),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1502 (
            .O(N__10903),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    InMux I__1501 (
            .O(N__10898),
            .I(N__10895));
    LocalMux I__1500 (
            .O(N__10895),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__1499 (
            .O(N__10892),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__1498 (
            .O(N__10889),
            .I(N__10882));
    InMux I__1497 (
            .O(N__10888),
            .I(N__10879));
    InMux I__1496 (
            .O(N__10887),
            .I(N__10874));
    InMux I__1495 (
            .O(N__10886),
            .I(N__10874));
    InMux I__1494 (
            .O(N__10885),
            .I(N__10871));
    LocalMux I__1493 (
            .O(N__10882),
            .I(N__10864));
    LocalMux I__1492 (
            .O(N__10879),
            .I(N__10864));
    LocalMux I__1491 (
            .O(N__10874),
            .I(N__10864));
    LocalMux I__1490 (
            .O(N__10871),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    Odrv12 I__1489 (
            .O(N__10864),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    CascadeMux I__1488 (
            .O(N__10859),
            .I(N__10856));
    InMux I__1487 (
            .O(N__10856),
            .I(N__10853));
    LocalMux I__1486 (
            .O(N__10853),
            .I(N__10850));
    Odrv12 I__1485 (
            .O(N__10850),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1484 (
            .O(N__10847),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    CascadeMux I__1483 (
            .O(N__10844),
            .I(N__10838));
    InMux I__1482 (
            .O(N__10843),
            .I(N__10834));
    InMux I__1481 (
            .O(N__10842),
            .I(N__10825));
    InMux I__1480 (
            .O(N__10841),
            .I(N__10825));
    InMux I__1479 (
            .O(N__10838),
            .I(N__10825));
    InMux I__1478 (
            .O(N__10837),
            .I(N__10825));
    LocalMux I__1477 (
            .O(N__10834),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1476 (
            .O(N__10825),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    CascadeMux I__1475 (
            .O(N__10820),
            .I(N__10817));
    InMux I__1474 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__1473 (
            .O(N__10814),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__1472 (
            .O(N__10811),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1471 (
            .O(N__10808),
            .I(N__10802));
    InMux I__1470 (
            .O(N__10807),
            .I(N__10802));
    LocalMux I__1469 (
            .O(N__10802),
            .I(N__10799));
    Span4Mux_h I__1468 (
            .O(N__10799),
            .I(N__10794));
    InMux I__1467 (
            .O(N__10798),
            .I(N__10791));
    InMux I__1466 (
            .O(N__10797),
            .I(N__10788));
    Odrv4 I__1465 (
            .O(N__10794),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1464 (
            .O(N__10791),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1463 (
            .O(N__10788),
            .I(\buart.Z_rx.N_27_0_i ));
    InMux I__1462 (
            .O(N__10781),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__1461 (
            .O(N__10778),
            .I(N__10775));
    InMux I__1460 (
            .O(N__10775),
            .I(N__10769));
    InMux I__1459 (
            .O(N__10774),
            .I(N__10762));
    InMux I__1458 (
            .O(N__10773),
            .I(N__10762));
    InMux I__1457 (
            .O(N__10772),
            .I(N__10762));
    LocalMux I__1456 (
            .O(N__10769),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1455 (
            .O(N__10762),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    InMux I__1454 (
            .O(N__10757),
            .I(N__10754));
    LocalMux I__1453 (
            .O(N__10754),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ));
    InMux I__1452 (
            .O(N__10751),
            .I(N__10747));
    InMux I__1451 (
            .O(N__10750),
            .I(N__10744));
    LocalMux I__1450 (
            .O(N__10747),
            .I(N__10741));
    LocalMux I__1449 (
            .O(N__10744),
            .I(N__10738));
    Odrv12 I__1448 (
            .O(N__10741),
            .I(\Lab_UT.di_ASones_0 ));
    Odrv4 I__1447 (
            .O(N__10738),
            .I(\Lab_UT.di_ASones_0 ));
    CEMux I__1446 (
            .O(N__10733),
            .I(N__10730));
    LocalMux I__1445 (
            .O(N__10730),
            .I(N__10727));
    Span4Mux_h I__1444 (
            .O(N__10727),
            .I(N__10724));
    Span4Mux_s0_h I__1443 (
            .O(N__10724),
            .I(N__10720));
    CEMux I__1442 (
            .O(N__10723),
            .I(N__10717));
    Odrv4 I__1441 (
            .O(N__10720),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    LocalMux I__1440 (
            .O(N__10717),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    CascadeMux I__1439 (
            .O(N__10712),
            .I(\buart.Z_rx.valid_0_cascade_ ));
    CascadeMux I__1438 (
            .O(N__10709),
            .I(\buart.Z_rx.idle_0_cascade_ ));
    CascadeMux I__1437 (
            .O(N__10706),
            .I(\buart.Z_rx.idle_cascade_ ));
    CascadeMux I__1436 (
            .O(N__10703),
            .I(\buart.Z_rx.N_27_0_i_cascade_ ));
    CascadeMux I__1435 (
            .O(N__10700),
            .I(\Lab_UT.three_2_1_cascade_ ));
    InMux I__1434 (
            .O(N__10697),
            .I(N__10694));
    LocalMux I__1433 (
            .O(N__10694),
            .I(\Lab_UT.didp.countrce3.q_5_2 ));
    CascadeMux I__1432 (
            .O(N__10691),
            .I(\Lab_UT.didp.countrce3.q_5_2_cascade_ ));
    CascadeMux I__1431 (
            .O(N__10688),
            .I(N__10684));
    InMux I__1430 (
            .O(N__10687),
            .I(N__10681));
    InMux I__1429 (
            .O(N__10684),
            .I(N__10678));
    LocalMux I__1428 (
            .O(N__10681),
            .I(\Lab_UT.didp.countrce3.q_fastZ0Z_2 ));
    LocalMux I__1427 (
            .O(N__10678),
            .I(\Lab_UT.didp.countrce3.q_fastZ0Z_2 ));
    InMux I__1426 (
            .O(N__10673),
            .I(N__10668));
    InMux I__1425 (
            .O(N__10672),
            .I(N__10665));
    InMux I__1424 (
            .O(N__10671),
            .I(N__10662));
    LocalMux I__1423 (
            .O(N__10668),
            .I(N__10659));
    LocalMux I__1422 (
            .O(N__10665),
            .I(\Lab_UT.di_AStens_2 ));
    LocalMux I__1421 (
            .O(N__10662),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__1420 (
            .O(N__10659),
            .I(\Lab_UT.di_AStens_2 ));
    CascadeMux I__1419 (
            .O(N__10652),
            .I(\Lab_UT.didp.did_alarmMatch_6_cascade_ ));
    InMux I__1418 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__1417 (
            .O(N__10646),
            .I(N__10643));
    Span4Mux_v I__1416 (
            .O(N__10643),
            .I(N__10640));
    Odrv4 I__1415 (
            .O(N__10640),
            .I(\Lab_UT.min2Z0Z_3 ));
    InMux I__1414 (
            .O(N__10637),
            .I(N__10634));
    LocalMux I__1413 (
            .O(N__10634),
            .I(N__10631));
    Odrv12 I__1412 (
            .O(N__10631),
            .I(\Lab_UT.min1Z0Z_1 ));
    InMux I__1411 (
            .O(N__10628),
            .I(N__10624));
    InMux I__1410 (
            .O(N__10627),
            .I(N__10621));
    LocalMux I__1409 (
            .O(N__10624),
            .I(N__10618));
    LocalMux I__1408 (
            .O(N__10621),
            .I(N__10615));
    Span4Mux_h I__1407 (
            .O(N__10618),
            .I(N__10612));
    Odrv4 I__1406 (
            .O(N__10615),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__1405 (
            .O(N__10612),
            .I(\Lab_UT.di_ASones_2 ));
    CascadeMux I__1404 (
            .O(N__10607),
            .I(N__10602));
    InMux I__1403 (
            .O(N__10606),
            .I(N__10589));
    InMux I__1402 (
            .O(N__10605),
            .I(N__10589));
    InMux I__1401 (
            .O(N__10602),
            .I(N__10586));
    InMux I__1400 (
            .O(N__10601),
            .I(N__10571));
    InMux I__1399 (
            .O(N__10600),
            .I(N__10571));
    InMux I__1398 (
            .O(N__10599),
            .I(N__10571));
    InMux I__1397 (
            .O(N__10598),
            .I(N__10571));
    InMux I__1396 (
            .O(N__10597),
            .I(N__10571));
    InMux I__1395 (
            .O(N__10596),
            .I(N__10571));
    InMux I__1394 (
            .O(N__10595),
            .I(N__10571));
    InMux I__1393 (
            .O(N__10594),
            .I(N__10564));
    LocalMux I__1392 (
            .O(N__10589),
            .I(N__10561));
    LocalMux I__1391 (
            .O(N__10586),
            .I(N__10558));
    LocalMux I__1390 (
            .O(N__10571),
            .I(N__10555));
    InMux I__1389 (
            .O(N__10570),
            .I(N__10548));
    InMux I__1388 (
            .O(N__10569),
            .I(N__10548));
    InMux I__1387 (
            .O(N__10568),
            .I(N__10548));
    CascadeMux I__1386 (
            .O(N__10567),
            .I(N__10545));
    LocalMux I__1385 (
            .O(N__10564),
            .I(N__10539));
    Span4Mux_v I__1384 (
            .O(N__10561),
            .I(N__10539));
    Span4Mux_v I__1383 (
            .O(N__10558),
            .I(N__10534));
    Span4Mux_s3_h I__1382 (
            .O(N__10555),
            .I(N__10534));
    LocalMux I__1381 (
            .O(N__10548),
            .I(N__10531));
    InMux I__1380 (
            .O(N__10545),
            .I(N__10526));
    InMux I__1379 (
            .O(N__10544),
            .I(N__10526));
    Odrv4 I__1378 (
            .O(N__10539),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1377 (
            .O(N__10534),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1376 (
            .O(N__10531),
            .I(vbuf_tx_data_rdy));
    LocalMux I__1375 (
            .O(N__10526),
            .I(vbuf_tx_data_rdy));
    InMux I__1374 (
            .O(N__10517),
            .I(N__10514));
    LocalMux I__1373 (
            .O(N__10514),
            .I(N__10510));
    CascadeMux I__1372 (
            .O(N__10513),
            .I(N__10507));
    Span4Mux_h I__1371 (
            .O(N__10510),
            .I(N__10502));
    InMux I__1370 (
            .O(N__10507),
            .I(N__10495));
    InMux I__1369 (
            .O(N__10506),
            .I(N__10495));
    InMux I__1368 (
            .O(N__10505),
            .I(N__10495));
    Odrv4 I__1367 (
            .O(N__10502),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__1366 (
            .O(N__10495),
            .I(\uu0.l_countZ0Z_10 ));
    InMux I__1365 (
            .O(N__10490),
            .I(N__10486));
    InMux I__1364 (
            .O(N__10489),
            .I(N__10481));
    LocalMux I__1363 (
            .O(N__10486),
            .I(N__10476));
    InMux I__1362 (
            .O(N__10485),
            .I(N__10471));
    InMux I__1361 (
            .O(N__10484),
            .I(N__10471));
    LocalMux I__1360 (
            .O(N__10481),
            .I(N__10468));
    InMux I__1359 (
            .O(N__10480),
            .I(N__10463));
    InMux I__1358 (
            .O(N__10479),
            .I(N__10463));
    Span4Mux_s1_h I__1357 (
            .O(N__10476),
            .I(N__10460));
    LocalMux I__1356 (
            .O(N__10471),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1355 (
            .O(N__10468),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1354 (
            .O(N__10463),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1353 (
            .O(N__10460),
            .I(\uu0.l_countZ0Z_8 ));
    InMux I__1352 (
            .O(N__10451),
            .I(N__10446));
    InMux I__1351 (
            .O(N__10450),
            .I(N__10441));
    InMux I__1350 (
            .O(N__10449),
            .I(N__10438));
    LocalMux I__1349 (
            .O(N__10446),
            .I(N__10435));
    InMux I__1348 (
            .O(N__10445),
            .I(N__10430));
    InMux I__1347 (
            .O(N__10444),
            .I(N__10430));
    LocalMux I__1346 (
            .O(N__10441),
            .I(N__10427));
    LocalMux I__1345 (
            .O(N__10438),
            .I(\uu0.l_countZ0Z_9 ));
    Odrv4 I__1344 (
            .O(N__10435),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1343 (
            .O(N__10430),
            .I(\uu0.l_countZ0Z_9 ));
    Odrv4 I__1342 (
            .O(N__10427),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__1341 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__1340 (
            .O(N__10415),
            .I(N__10412));
    Odrv4 I__1339 (
            .O(N__10412),
            .I(\uu0.un143_ci_0 ));
    CEMux I__1338 (
            .O(N__10409),
            .I(N__10406));
    LocalMux I__1337 (
            .O(N__10406),
            .I(N__10402));
    CEMux I__1336 (
            .O(N__10405),
            .I(N__10399));
    Span4Mux_v I__1335 (
            .O(N__10402),
            .I(N__10394));
    LocalMux I__1334 (
            .O(N__10399),
            .I(N__10394));
    Span4Mux_v I__1333 (
            .O(N__10394),
            .I(N__10391));
    Span4Mux_s2_h I__1332 (
            .O(N__10391),
            .I(N__10388));
    Odrv4 I__1331 (
            .O(N__10388),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    CascadeMux I__1330 (
            .O(N__10385),
            .I(N__10382));
    InMux I__1329 (
            .O(N__10382),
            .I(N__10379));
    LocalMux I__1328 (
            .O(N__10379),
            .I(N__10376));
    Odrv12 I__1327 (
            .O(N__10376),
            .I(\resetGen.reset_count_2_0_4 ));
    InMux I__1326 (
            .O(N__10373),
            .I(N__10370));
    LocalMux I__1325 (
            .O(N__10370),
            .I(\Lab_UT.dispString.N_46 ));
    CascadeMux I__1324 (
            .O(N__10367),
            .I(N__10364));
    InMux I__1323 (
            .O(N__10364),
            .I(N__10361));
    LocalMux I__1322 (
            .O(N__10361),
            .I(\Lab_UT.min2Z0Z_1 ));
    InMux I__1321 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__1320 (
            .O(N__10355),
            .I(\Lab_UT.min2Z0Z_2 ));
    CascadeMux I__1319 (
            .O(N__10352),
            .I(N__10349));
    InMux I__1318 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__1317 (
            .O(N__10346),
            .I(\Lab_UT.sec1Z0Z_2 ));
    CascadeMux I__1316 (
            .O(N__10343),
            .I(\Lab_UT.dicLdAStens_0_cascade_ ));
    InMux I__1315 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__1314 (
            .O(N__10337),
            .I(\Lab_UT.alarmcharZ0Z_5 ));
    CascadeMux I__1313 (
            .O(N__10334),
            .I(\Lab_UT.dispString.m35_ns_1_cascade_ ));
    InMux I__1312 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__1311 (
            .O(N__10328),
            .I(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ));
    CascadeMux I__1310 (
            .O(N__10325),
            .I(N__10322));
    InMux I__1309 (
            .O(N__10322),
            .I(N__10319));
    LocalMux I__1308 (
            .O(N__10319),
            .I(\Lab_UT.sec2Z0Z_0 ));
    InMux I__1307 (
            .O(N__10316),
            .I(N__10313));
    LocalMux I__1306 (
            .O(N__10313),
            .I(\Lab_UT.alarmcharZ0Z_0 ));
    CascadeMux I__1305 (
            .O(N__10310),
            .I(\Lab_UT.dispString.m32_ns_1_cascade_ ));
    CascadeMux I__1304 (
            .O(N__10307),
            .I(N__10304));
    InMux I__1303 (
            .O(N__10304),
            .I(N__10301));
    LocalMux I__1302 (
            .O(N__10301),
            .I(\Lab_UT.sec1Z0Z_3 ));
    CascadeMux I__1301 (
            .O(N__10298),
            .I(N__10295));
    InMux I__1300 (
            .O(N__10295),
            .I(N__10292));
    LocalMux I__1299 (
            .O(N__10292),
            .I(\Lab_UT.sec2Z0Z_1 ));
    CascadeMux I__1298 (
            .O(N__10289),
            .I(\Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ));
    CEMux I__1297 (
            .O(N__10286),
            .I(N__10281));
    CEMux I__1296 (
            .O(N__10285),
            .I(N__10278));
    CEMux I__1295 (
            .O(N__10284),
            .I(N__10275));
    LocalMux I__1294 (
            .O(N__10281),
            .I(N__10270));
    LocalMux I__1293 (
            .O(N__10278),
            .I(N__10270));
    LocalMux I__1292 (
            .O(N__10275),
            .I(N__10267));
    Span4Mux_v I__1291 (
            .O(N__10270),
            .I(N__10264));
    Span4Mux_h I__1290 (
            .O(N__10267),
            .I(N__10261));
    Odrv4 I__1289 (
            .O(N__10264),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__1288 (
            .O(N__10261),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1287 (
            .O(N__10256),
            .I(N__10253));
    LocalMux I__1286 (
            .O(N__10253),
            .I(N__10250));
    Span4Mux_h I__1285 (
            .O(N__10250),
            .I(N__10246));
    InMux I__1284 (
            .O(N__10249),
            .I(N__10243));
    Odrv4 I__1283 (
            .O(N__10246),
            .I(\uu2.un1_l_count_1_0 ));
    LocalMux I__1282 (
            .O(N__10243),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1281 (
            .O(N__10238),
            .I(N__10235));
    LocalMux I__1280 (
            .O(N__10235),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1279 (
            .O(N__10232),
            .I(N__10229));
    LocalMux I__1278 (
            .O(N__10229),
            .I(\uu2.mem0.w_data_0 ));
    InMux I__1277 (
            .O(N__10226),
            .I(N__10223));
    LocalMux I__1276 (
            .O(N__10223),
            .I(\uu2.mem0.N_30_i_0 ));
    CascadeMux I__1275 (
            .O(N__10220),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_ ));
    InMux I__1274 (
            .O(N__10217),
            .I(N__10214));
    LocalMux I__1273 (
            .O(N__10214),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1272 (
            .O(N__10211),
            .I(N__10207));
    InMux I__1271 (
            .O(N__10210),
            .I(N__10204));
    LocalMux I__1270 (
            .O(N__10207),
            .I(N__10198));
    LocalMux I__1269 (
            .O(N__10204),
            .I(N__10198));
    CascadeMux I__1268 (
            .O(N__10203),
            .I(N__10194));
    Span4Mux_v I__1267 (
            .O(N__10198),
            .I(N__10190));
    InMux I__1266 (
            .O(N__10197),
            .I(N__10183));
    InMux I__1265 (
            .O(N__10194),
            .I(N__10183));
    InMux I__1264 (
            .O(N__10193),
            .I(N__10183));
    Odrv4 I__1263 (
            .O(N__10190),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__1262 (
            .O(N__10183),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__1261 (
            .O(N__10178),
            .I(\uu2.vbuf_raddr.un448_ci_0_cascade_ ));
    CascadeMux I__1260 (
            .O(N__10175),
            .I(N__10172));
    InMux I__1259 (
            .O(N__10172),
            .I(N__10168));
    InMux I__1258 (
            .O(N__10171),
            .I(N__10165));
    LocalMux I__1257 (
            .O(N__10168),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1256 (
            .O(N__10165),
            .I(\uu2.r_addrZ0Z_8 ));
    InMux I__1255 (
            .O(N__10160),
            .I(N__10157));
    LocalMux I__1254 (
            .O(N__10157),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__1253 (
            .O(N__10154),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1252 (
            .O(N__10151),
            .I(N__10148));
    InMux I__1251 (
            .O(N__10148),
            .I(N__10143));
    InMux I__1250 (
            .O(N__10147),
            .I(N__10138));
    InMux I__1249 (
            .O(N__10146),
            .I(N__10138));
    LocalMux I__1248 (
            .O(N__10143),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1247 (
            .O(N__10138),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__1246 (
            .O(N__10133),
            .I(N__10127));
    InMux I__1245 (
            .O(N__10132),
            .I(N__10127));
    LocalMux I__1244 (
            .O(N__10127),
            .I(N__10122));
    InMux I__1243 (
            .O(N__10126),
            .I(N__10117));
    InMux I__1242 (
            .O(N__10125),
            .I(N__10117));
    Odrv4 I__1241 (
            .O(N__10122),
            .I(\uu2.un404_ci_0 ));
    LocalMux I__1240 (
            .O(N__10117),
            .I(\uu2.un404_ci_0 ));
    CascadeMux I__1239 (
            .O(N__10112),
            .I(N__10105));
    InMux I__1238 (
            .O(N__10111),
            .I(N__10100));
    InMux I__1237 (
            .O(N__10110),
            .I(N__10100));
    InMux I__1236 (
            .O(N__10109),
            .I(N__10095));
    InMux I__1235 (
            .O(N__10108),
            .I(N__10095));
    InMux I__1234 (
            .O(N__10105),
            .I(N__10092));
    LocalMux I__1233 (
            .O(N__10100),
            .I(N__10087));
    LocalMux I__1232 (
            .O(N__10095),
            .I(N__10087));
    LocalMux I__1231 (
            .O(N__10092),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1230 (
            .O(N__10087),
            .I(\uu2.r_addrZ0Z_4 ));
    CascadeMux I__1229 (
            .O(N__10082),
            .I(\uu2.un404_ci_0_cascade_ ));
    CascadeMux I__1228 (
            .O(N__10079),
            .I(N__10073));
    CascadeMux I__1227 (
            .O(N__10078),
            .I(N__10070));
    InMux I__1226 (
            .O(N__10077),
            .I(N__10067));
    InMux I__1225 (
            .O(N__10076),
            .I(N__10064));
    InMux I__1224 (
            .O(N__10073),
            .I(N__10061));
    InMux I__1223 (
            .O(N__10070),
            .I(N__10058));
    LocalMux I__1222 (
            .O(N__10067),
            .I(N__10053));
    LocalMux I__1221 (
            .O(N__10064),
            .I(N__10053));
    LocalMux I__1220 (
            .O(N__10061),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1219 (
            .O(N__10058),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__1218 (
            .O(N__10053),
            .I(\uu2.r_addrZ0Z_5 ));
    CascadeMux I__1217 (
            .O(N__10046),
            .I(N__10043));
    InMux I__1216 (
            .O(N__10043),
            .I(N__10037));
    InMux I__1215 (
            .O(N__10042),
            .I(N__10032));
    InMux I__1214 (
            .O(N__10041),
            .I(N__10032));
    InMux I__1213 (
            .O(N__10040),
            .I(N__10029));
    LocalMux I__1212 (
            .O(N__10037),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1211 (
            .O(N__10032),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1210 (
            .O(N__10029),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1209 (
            .O(N__10022),
            .I(N__10019));
    InMux I__1208 (
            .O(N__10019),
            .I(N__10016));
    LocalMux I__1207 (
            .O(N__10016),
            .I(N__10012));
    CascadeMux I__1206 (
            .O(N__10015),
            .I(N__10009));
    Span4Mux_v I__1205 (
            .O(N__10012),
            .I(N__10004));
    InMux I__1204 (
            .O(N__10009),
            .I(N__10001));
    InMux I__1203 (
            .O(N__10008),
            .I(N__9996));
    InMux I__1202 (
            .O(N__10007),
            .I(N__9996));
    Odrv4 I__1201 (
            .O(N__10004),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1200 (
            .O(N__10001),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1199 (
            .O(N__9996),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1198 (
            .O(N__9989),
            .I(N__9986));
    InMux I__1197 (
            .O(N__9986),
            .I(N__9983));
    LocalMux I__1196 (
            .O(N__9983),
            .I(N__9976));
    InMux I__1195 (
            .O(N__9982),
            .I(N__9971));
    InMux I__1194 (
            .O(N__9981),
            .I(N__9971));
    InMux I__1193 (
            .O(N__9980),
            .I(N__9966));
    InMux I__1192 (
            .O(N__9979),
            .I(N__9966));
    Odrv4 I__1191 (
            .O(N__9976),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1190 (
            .O(N__9971),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1189 (
            .O(N__9966),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1188 (
            .O(N__9959),
            .I(N__9956));
    InMux I__1187 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__1186 (
            .O(N__9953),
            .I(N__9950));
    Span4Mux_s3_h I__1185 (
            .O(N__9950),
            .I(N__9942));
    InMux I__1184 (
            .O(N__9949),
            .I(N__9935));
    InMux I__1183 (
            .O(N__9948),
            .I(N__9935));
    InMux I__1182 (
            .O(N__9947),
            .I(N__9935));
    InMux I__1181 (
            .O(N__9946),
            .I(N__9930));
    InMux I__1180 (
            .O(N__9945),
            .I(N__9930));
    Odrv4 I__1179 (
            .O(N__9942),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1178 (
            .O(N__9935),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1177 (
            .O(N__9930),
            .I(\uu2.r_addrZ0Z_0 ));
    CascadeMux I__1176 (
            .O(N__9923),
            .I(N__9918));
    CascadeMux I__1175 (
            .O(N__9922),
            .I(N__9915));
    CascadeMux I__1174 (
            .O(N__9921),
            .I(N__9912));
    InMux I__1173 (
            .O(N__9918),
            .I(N__9909));
    InMux I__1172 (
            .O(N__9915),
            .I(N__9904));
    InMux I__1171 (
            .O(N__9912),
            .I(N__9904));
    LocalMux I__1170 (
            .O(N__9909),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1169 (
            .O(N__9904),
            .I(\uu2.r_addrZ0Z_3 ));
    CEMux I__1168 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__1167 (
            .O(N__9896),
            .I(N__9893));
    Span4Mux_v I__1166 (
            .O(N__9893),
            .I(N__9890));
    Odrv4 I__1165 (
            .O(N__9890),
            .I(\uu2.trig_rd_is_det_0 ));
    InMux I__1164 (
            .O(N__9887),
            .I(N__9882));
    InMux I__1163 (
            .O(N__9886),
            .I(N__9879));
    CascadeMux I__1162 (
            .O(N__9885),
            .I(N__9875));
    LocalMux I__1161 (
            .O(N__9882),
            .I(N__9870));
    LocalMux I__1160 (
            .O(N__9879),
            .I(N__9870));
    InMux I__1159 (
            .O(N__9878),
            .I(N__9865));
    InMux I__1158 (
            .O(N__9875),
            .I(N__9865));
    Odrv4 I__1157 (
            .O(N__9870),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__1156 (
            .O(N__9865),
            .I(\uu0.un154_ci_9 ));
    InMux I__1155 (
            .O(N__9860),
            .I(N__9851));
    InMux I__1154 (
            .O(N__9859),
            .I(N__9851));
    InMux I__1153 (
            .O(N__9858),
            .I(N__9851));
    LocalMux I__1152 (
            .O(N__9851),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__1151 (
            .O(N__9848),
            .I(N__9845));
    LocalMux I__1150 (
            .O(N__9845),
            .I(N__9842));
    Odrv12 I__1149 (
            .O(N__9842),
            .I(\uu0.un165_ci_0 ));
    InMux I__1148 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__1147 (
            .O(N__9836),
            .I(N__9833));
    Odrv4 I__1146 (
            .O(N__9833),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1145 (
            .O(N__9830),
            .I(N__9827));
    LocalMux I__1144 (
            .O(N__9827),
            .I(N__9823));
    InMux I__1143 (
            .O(N__9826),
            .I(N__9820));
    Span4Mux_h I__1142 (
            .O(N__9823),
            .I(N__9817));
    LocalMux I__1141 (
            .O(N__9820),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    Odrv4 I__1140 (
            .O(N__9817),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    CascadeMux I__1139 (
            .O(N__9812),
            .I(\uu2.trig_rd_is_det_cascade_ ));
    CascadeMux I__1138 (
            .O(N__9809),
            .I(N__9804));
    CascadeMux I__1137 (
            .O(N__9808),
            .I(N__9801));
    InMux I__1136 (
            .O(N__9807),
            .I(N__9798));
    InMux I__1135 (
            .O(N__9804),
            .I(N__9795));
    InMux I__1134 (
            .O(N__9801),
            .I(N__9792));
    LocalMux I__1133 (
            .O(N__9798),
            .I(N__9789));
    LocalMux I__1132 (
            .O(N__9795),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__1131 (
            .O(N__9792),
            .I(\uu0.l_countZ0Z_11 ));
    Odrv4 I__1130 (
            .O(N__9789),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__1129 (
            .O(N__9782),
            .I(N__9779));
    InMux I__1128 (
            .O(N__9779),
            .I(N__9773));
    InMux I__1127 (
            .O(N__9778),
            .I(N__9770));
    InMux I__1126 (
            .O(N__9777),
            .I(N__9765));
    InMux I__1125 (
            .O(N__9776),
            .I(N__9765));
    LocalMux I__1124 (
            .O(N__9773),
            .I(N__9762));
    LocalMux I__1123 (
            .O(N__9770),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__1122 (
            .O(N__9765),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1121 (
            .O(N__9762),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__1120 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__1119 (
            .O(N__9752),
            .I(\uu0.un4_l_count_11 ));
    InMux I__1118 (
            .O(N__9749),
            .I(N__9746));
    LocalMux I__1117 (
            .O(N__9746),
            .I(\uu0.un4_l_count_16 ));
    CascadeMux I__1116 (
            .O(N__9743),
            .I(N__9740));
    InMux I__1115 (
            .O(N__9740),
            .I(N__9730));
    InMux I__1114 (
            .O(N__9739),
            .I(N__9730));
    InMux I__1113 (
            .O(N__9738),
            .I(N__9730));
    InMux I__1112 (
            .O(N__9737),
            .I(N__9727));
    LocalMux I__1111 (
            .O(N__9730),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1110 (
            .O(N__9727),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__1109 (
            .O(N__9722),
            .I(N__9717));
    CascadeMux I__1108 (
            .O(N__9721),
            .I(N__9714));
    InMux I__1107 (
            .O(N__9720),
            .I(N__9707));
    InMux I__1106 (
            .O(N__9717),
            .I(N__9707));
    InMux I__1105 (
            .O(N__9714),
            .I(N__9707));
    LocalMux I__1104 (
            .O(N__9707),
            .I(N__9704));
    Odrv4 I__1103 (
            .O(N__9704),
            .I(\uu0.un198_ci_2 ));
    CascadeMux I__1102 (
            .O(N__9701),
            .I(N__9696));
    InMux I__1101 (
            .O(N__9700),
            .I(N__9691));
    InMux I__1100 (
            .O(N__9699),
            .I(N__9691));
    InMux I__1099 (
            .O(N__9696),
            .I(N__9688));
    LocalMux I__1098 (
            .O(N__9691),
            .I(\uu0.l_countZ0Z_17 ));
    LocalMux I__1097 (
            .O(N__9688),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__1096 (
            .O(N__9683),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__1095 (
            .O(N__9680),
            .I(N__9676));
    InMux I__1094 (
            .O(N__9679),
            .I(N__9673));
    LocalMux I__1093 (
            .O(N__9676),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__1092 (
            .O(N__9673),
            .I(\uu0.l_countZ0Z_18 ));
    CascadeMux I__1091 (
            .O(N__9668),
            .I(N__9664));
    InMux I__1090 (
            .O(N__9667),
            .I(N__9661));
    InMux I__1089 (
            .O(N__9664),
            .I(N__9658));
    LocalMux I__1088 (
            .O(N__9661),
            .I(N__9655));
    LocalMux I__1087 (
            .O(N__9658),
            .I(\uu0.l_countZ0Z_13 ));
    Odrv4 I__1086 (
            .O(N__9655),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__1085 (
            .O(N__9650),
            .I(N__9641));
    InMux I__1084 (
            .O(N__9649),
            .I(N__9641));
    InMux I__1083 (
            .O(N__9648),
            .I(N__9641));
    LocalMux I__1082 (
            .O(N__9641),
            .I(N__9637));
    InMux I__1081 (
            .O(N__9640),
            .I(N__9634));
    Odrv4 I__1080 (
            .O(N__9637),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__1079 (
            .O(N__9634),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__1078 (
            .O(N__9629),
            .I(N__9624));
    InMux I__1077 (
            .O(N__9628),
            .I(N__9607));
    InMux I__1076 (
            .O(N__9627),
            .I(N__9607));
    InMux I__1075 (
            .O(N__9624),
            .I(N__9607));
    InMux I__1074 (
            .O(N__9623),
            .I(N__9607));
    InMux I__1073 (
            .O(N__9622),
            .I(N__9602));
    InMux I__1072 (
            .O(N__9621),
            .I(N__9602));
    InMux I__1071 (
            .O(N__9620),
            .I(N__9599));
    InMux I__1070 (
            .O(N__9619),
            .I(N__9590));
    InMux I__1069 (
            .O(N__9618),
            .I(N__9590));
    InMux I__1068 (
            .O(N__9617),
            .I(N__9590));
    InMux I__1067 (
            .O(N__9616),
            .I(N__9590));
    LocalMux I__1066 (
            .O(N__9607),
            .I(N__9587));
    LocalMux I__1065 (
            .O(N__9602),
            .I(\uu0.un110_ci ));
    LocalMux I__1064 (
            .O(N__9599),
            .I(\uu0.un110_ci ));
    LocalMux I__1063 (
            .O(N__9590),
            .I(\uu0.un110_ci ));
    Odrv4 I__1062 (
            .O(N__9587),
            .I(\uu0.un110_ci ));
    InMux I__1061 (
            .O(N__9578),
            .I(N__9572));
    InMux I__1060 (
            .O(N__9577),
            .I(N__9562));
    InMux I__1059 (
            .O(N__9576),
            .I(N__9562));
    InMux I__1058 (
            .O(N__9575),
            .I(N__9562));
    LocalMux I__1057 (
            .O(N__9572),
            .I(N__9553));
    InMux I__1056 (
            .O(N__9571),
            .I(N__9546));
    InMux I__1055 (
            .O(N__9570),
            .I(N__9546));
    InMux I__1054 (
            .O(N__9569),
            .I(N__9546));
    LocalMux I__1053 (
            .O(N__9562),
            .I(N__9543));
    InMux I__1052 (
            .O(N__9561),
            .I(N__9538));
    InMux I__1051 (
            .O(N__9560),
            .I(N__9538));
    InMux I__1050 (
            .O(N__9559),
            .I(N__9531));
    InMux I__1049 (
            .O(N__9558),
            .I(N__9531));
    InMux I__1048 (
            .O(N__9557),
            .I(N__9531));
    InMux I__1047 (
            .O(N__9556),
            .I(N__9528));
    Odrv12 I__1046 (
            .O(N__9553),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1045 (
            .O(N__9546),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1044 (
            .O(N__9543),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1043 (
            .O(N__9538),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1042 (
            .O(N__9531),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1041 (
            .O(N__9528),
            .I(\uu0.un4_l_count_0 ));
    CEMux I__1040 (
            .O(N__9515),
            .I(N__9503));
    CEMux I__1039 (
            .O(N__9514),
            .I(N__9503));
    CEMux I__1038 (
            .O(N__9513),
            .I(N__9503));
    CEMux I__1037 (
            .O(N__9512),
            .I(N__9503));
    GlobalMux I__1036 (
            .O(N__9503),
            .I(N__9500));
    gio2CtrlBuf I__1035 (
            .O(N__9500),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__1034 (
            .O(N__9497),
            .I(\uu0.un154_ci_9_cascade_ ));
    InMux I__1033 (
            .O(N__9494),
            .I(N__9486));
    InMux I__1032 (
            .O(N__9493),
            .I(N__9486));
    InMux I__1031 (
            .O(N__9492),
            .I(N__9483));
    InMux I__1030 (
            .O(N__9491),
            .I(N__9480));
    LocalMux I__1029 (
            .O(N__9486),
            .I(\uu0.un66_ci ));
    LocalMux I__1028 (
            .O(N__9483),
            .I(\uu0.un66_ci ));
    LocalMux I__1027 (
            .O(N__9480),
            .I(\uu0.un66_ci ));
    InMux I__1026 (
            .O(N__9473),
            .I(N__9461));
    InMux I__1025 (
            .O(N__9472),
            .I(N__9461));
    InMux I__1024 (
            .O(N__9471),
            .I(N__9461));
    InMux I__1023 (
            .O(N__9470),
            .I(N__9461));
    LocalMux I__1022 (
            .O(N__9461),
            .I(\uu0.l_countZ0Z_14 ));
    CascadeMux I__1021 (
            .O(N__9458),
            .I(N__9453));
    InMux I__1020 (
            .O(N__9457),
            .I(N__9448));
    InMux I__1019 (
            .O(N__9456),
            .I(N__9448));
    InMux I__1018 (
            .O(N__9453),
            .I(N__9445));
    LocalMux I__1017 (
            .O(N__9448),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__1016 (
            .O(N__9445),
            .I(\uu0.l_countZ0Z_15 ));
    InMux I__1015 (
            .O(N__9440),
            .I(N__9434));
    InMux I__1014 (
            .O(N__9439),
            .I(N__9431));
    InMux I__1013 (
            .O(N__9438),
            .I(N__9426));
    InMux I__1012 (
            .O(N__9437),
            .I(N__9426));
    LocalMux I__1011 (
            .O(N__9434),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__1010 (
            .O(N__9431),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__1009 (
            .O(N__9426),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__1008 (
            .O(N__9419),
            .I(N__9414));
    InMux I__1007 (
            .O(N__9418),
            .I(N__9411));
    InMux I__1006 (
            .O(N__9417),
            .I(N__9408));
    LocalMux I__1005 (
            .O(N__9414),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__1004 (
            .O(N__9411),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__1003 (
            .O(N__9408),
            .I(\uu0.l_countZ0Z_7 ));
    InMux I__1002 (
            .O(N__9401),
            .I(N__9394));
    InMux I__1001 (
            .O(N__9400),
            .I(N__9394));
    InMux I__1000 (
            .O(N__9399),
            .I(N__9391));
    LocalMux I__999 (
            .O(N__9394),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__998 (
            .O(N__9391),
            .I(\uu0.l_countZ0Z_3 ));
    InMux I__997 (
            .O(N__9386),
            .I(N__9383));
    LocalMux I__996 (
            .O(N__9383),
            .I(\uu0.un4_l_count_14 ));
    CascadeMux I__995 (
            .O(N__9380),
            .I(N__9377));
    InMux I__994 (
            .O(N__9377),
            .I(N__9364));
    InMux I__993 (
            .O(N__9376),
            .I(N__9364));
    InMux I__992 (
            .O(N__9375),
            .I(N__9364));
    InMux I__991 (
            .O(N__9374),
            .I(N__9364));
    CascadeMux I__990 (
            .O(N__9373),
            .I(N__9360));
    LocalMux I__989 (
            .O(N__9364),
            .I(N__9357));
    InMux I__988 (
            .O(N__9363),
            .I(N__9354));
    InMux I__987 (
            .O(N__9360),
            .I(N__9351));
    Odrv4 I__986 (
            .O(N__9357),
            .I(\uu0.l_precountZ0Z_0 ));
    LocalMux I__985 (
            .O(N__9354),
            .I(\uu0.l_precountZ0Z_0 ));
    LocalMux I__984 (
            .O(N__9351),
            .I(\uu0.l_precountZ0Z_0 ));
    InMux I__983 (
            .O(N__9344),
            .I(N__9341));
    LocalMux I__982 (
            .O(N__9341),
            .I(\uu0.un4_l_count_13 ));
    InMux I__981 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__980 (
            .O(N__9335),
            .I(\uu0.un4_l_count_12 ));
    CascadeMux I__979 (
            .O(N__9332),
            .I(\uu0.un4_l_count_18_cascade_ ));
    InMux I__978 (
            .O(N__9329),
            .I(N__9326));
    LocalMux I__977 (
            .O(N__9326),
            .I(N__9323));
    Odrv4 I__976 (
            .O(N__9323),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__975 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__974 (
            .O(N__9317),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__973 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__972 (
            .O(N__9311),
            .I(N__9308));
    Span4Mux_s0_h I__971 (
            .O(N__9308),
            .I(N__9305));
    Span4Mux_v I__970 (
            .O(N__9305),
            .I(N__9302));
    Odrv4 I__969 (
            .O(N__9302),
            .I(o_serial_data_c));
    CascadeMux I__968 (
            .O(N__9299),
            .I(N__9296));
    InMux I__967 (
            .O(N__9296),
            .I(N__9292));
    InMux I__966 (
            .O(N__9295),
            .I(N__9289));
    LocalMux I__965 (
            .O(N__9292),
            .I(\uu0.un88_ci_3 ));
    LocalMux I__964 (
            .O(N__9289),
            .I(\uu0.un88_ci_3 ));
    InMux I__963 (
            .O(N__9284),
            .I(N__9279));
    InMux I__962 (
            .O(N__9283),
            .I(N__9276));
    InMux I__961 (
            .O(N__9282),
            .I(N__9273));
    LocalMux I__960 (
            .O(N__9279),
            .I(N__9270));
    LocalMux I__959 (
            .O(N__9276),
            .I(\uu0.l_countZ0Z_5 ));
    LocalMux I__958 (
            .O(N__9273),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv4 I__957 (
            .O(N__9270),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__956 (
            .O(N__9263),
            .I(\uu0.un187_ci_1_cascade_ ));
    InMux I__955 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__954 (
            .O(N__9257),
            .I(vbuf_tx_data_0));
    InMux I__953 (
            .O(N__9254),
            .I(N__9251));
    LocalMux I__952 (
            .O(N__9251),
            .I(vbuf_tx_data_7));
    InMux I__951 (
            .O(N__9248),
            .I(N__9245));
    LocalMux I__950 (
            .O(N__9245),
            .I(N__9242));
    Odrv4 I__949 (
            .O(N__9242),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    InMux I__948 (
            .O(N__9239),
            .I(N__9236));
    LocalMux I__947 (
            .O(N__9236),
            .I(vbuf_tx_data_1));
    InMux I__946 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__945 (
            .O(N__9230),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__944 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__943 (
            .O(N__9224),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__942 (
            .O(N__9221),
            .I(N__9218));
    LocalMux I__941 (
            .O(N__9218),
            .I(vbuf_tx_data_3));
    InMux I__940 (
            .O(N__9215),
            .I(N__9212));
    LocalMux I__939 (
            .O(N__9212),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__938 (
            .O(N__9209),
            .I(N__9206));
    LocalMux I__937 (
            .O(N__9206),
            .I(vbuf_tx_data_4));
    InMux I__936 (
            .O(N__9203),
            .I(N__9200));
    LocalMux I__935 (
            .O(N__9200),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__934 (
            .O(N__9197),
            .I(N__9194));
    LocalMux I__933 (
            .O(N__9194),
            .I(N__9191));
    Odrv4 I__932 (
            .O(N__9191),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__931 (
            .O(N__9188),
            .I(N__9185));
    LocalMux I__930 (
            .O(N__9185),
            .I(vbuf_tx_data_5));
    InMux I__929 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__928 (
            .O(N__9179),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__927 (
            .O(N__9176),
            .I(N__9173));
    LocalMux I__926 (
            .O(N__9173),
            .I(N__9170));
    Span12Mux_s2_h I__925 (
            .O(N__9170),
            .I(N__9167));
    Odrv12 I__924 (
            .O(N__9167),
            .I(\uu2.r_data_wire_2 ));
    InMux I__923 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__922 (
            .O(N__9161),
            .I(vbuf_tx_data_2));
    InMux I__921 (
            .O(N__9158),
            .I(N__9151));
    InMux I__920 (
            .O(N__9157),
            .I(N__9148));
    InMux I__919 (
            .O(N__9156),
            .I(N__9141));
    InMux I__918 (
            .O(N__9155),
            .I(N__9141));
    InMux I__917 (
            .O(N__9154),
            .I(N__9141));
    LocalMux I__916 (
            .O(N__9151),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__915 (
            .O(N__9148),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__914 (
            .O(N__9141),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__913 (
            .O(N__9134),
            .I(N__9129));
    InMux I__912 (
            .O(N__9133),
            .I(N__9123));
    InMux I__911 (
            .O(N__9132),
            .I(N__9120));
    LocalMux I__910 (
            .O(N__9129),
            .I(N__9117));
    InMux I__909 (
            .O(N__9128),
            .I(N__9114));
    InMux I__908 (
            .O(N__9127),
            .I(N__9109));
    InMux I__907 (
            .O(N__9126),
            .I(N__9109));
    LocalMux I__906 (
            .O(N__9123),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__905 (
            .O(N__9120),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__904 (
            .O(N__9117),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__903 (
            .O(N__9114),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__902 (
            .O(N__9109),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__901 (
            .O(N__9098),
            .I(N__9092));
    InMux I__900 (
            .O(N__9097),
            .I(N__9092));
    LocalMux I__899 (
            .O(N__9092),
            .I(\uu2.un284_ci ));
    InMux I__898 (
            .O(N__9089),
            .I(N__9086));
    LocalMux I__897 (
            .O(N__9086),
            .I(N__9083));
    Odrv4 I__896 (
            .O(N__9083),
            .I(\uu2.r_data_wire_0 ));
    InMux I__895 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__894 (
            .O(N__9077),
            .I(N__9074));
    Odrv4 I__893 (
            .O(N__9074),
            .I(\uu2.r_data_wire_1 ));
    InMux I__892 (
            .O(N__9071),
            .I(N__9068));
    LocalMux I__891 (
            .O(N__9068),
            .I(N__9065));
    Odrv4 I__890 (
            .O(N__9065),
            .I(\uu2.r_data_wire_3 ));
    InMux I__889 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__888 (
            .O(N__9059),
            .I(\uu2.r_data_wire_4 ));
    InMux I__887 (
            .O(N__9056),
            .I(N__9053));
    LocalMux I__886 (
            .O(N__9053),
            .I(\uu2.r_data_wire_5 ));
    InMux I__885 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__884 (
            .O(N__9047),
            .I(\uu2.r_data_wire_6 ));
    InMux I__883 (
            .O(N__9044),
            .I(N__9041));
    LocalMux I__882 (
            .O(N__9041),
            .I(N__9038));
    Odrv4 I__881 (
            .O(N__9038),
            .I(vbuf_tx_data_6));
    InMux I__880 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__879 (
            .O(N__9032),
            .I(\uu2.r_data_wire_7 ));
    InMux I__878 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__877 (
            .O(N__9026),
            .I(N__9023));
    IoSpan4Mux I__876 (
            .O(N__9023),
            .I(N__9020));
    Odrv4 I__875 (
            .O(N__9020),
            .I(uart_RXD));
    InMux I__874 (
            .O(N__9017),
            .I(N__9010));
    InMux I__873 (
            .O(N__9016),
            .I(N__9007));
    InMux I__872 (
            .O(N__9015),
            .I(N__9000));
    InMux I__871 (
            .O(N__9014),
            .I(N__9000));
    InMux I__870 (
            .O(N__9013),
            .I(N__9000));
    LocalMux I__869 (
            .O(N__9010),
            .I(\uu2.un306_ci ));
    LocalMux I__868 (
            .O(N__9007),
            .I(\uu2.un306_ci ));
    LocalMux I__867 (
            .O(N__9000),
            .I(\uu2.un306_ci ));
    CascadeMux I__866 (
            .O(N__8993),
            .I(N__8987));
    InMux I__865 (
            .O(N__8992),
            .I(N__8983));
    InMux I__864 (
            .O(N__8991),
            .I(N__8980));
    InMux I__863 (
            .O(N__8990),
            .I(N__8977));
    InMux I__862 (
            .O(N__8987),
            .I(N__8972));
    InMux I__861 (
            .O(N__8986),
            .I(N__8972));
    LocalMux I__860 (
            .O(N__8983),
            .I(N__8969));
    LocalMux I__859 (
            .O(N__8980),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__858 (
            .O(N__8977),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__857 (
            .O(N__8972),
            .I(\uu2.l_countZ0Z_4 ));
    Odrv4 I__856 (
            .O(N__8969),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__855 (
            .O(N__8960),
            .I(N__8955));
    InMux I__854 (
            .O(N__8959),
            .I(N__8952));
    InMux I__853 (
            .O(N__8958),
            .I(N__8949));
    LocalMux I__852 (
            .O(N__8955),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__851 (
            .O(N__8952),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__850 (
            .O(N__8949),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__849 (
            .O(N__8942),
            .I(N__8937));
    InMux I__848 (
            .O(N__8941),
            .I(N__8934));
    InMux I__847 (
            .O(N__8940),
            .I(N__8931));
    LocalMux I__846 (
            .O(N__8937),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__845 (
            .O(N__8934),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__844 (
            .O(N__8931),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__843 (
            .O(N__8924),
            .I(N__8919));
    CascadeMux I__842 (
            .O(N__8923),
            .I(N__8916));
    InMux I__841 (
            .O(N__8922),
            .I(N__8909));
    InMux I__840 (
            .O(N__8919),
            .I(N__8909));
    InMux I__839 (
            .O(N__8916),
            .I(N__8909));
    LocalMux I__838 (
            .O(N__8909),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__837 (
            .O(N__8906),
            .I(N__8900));
    InMux I__836 (
            .O(N__8905),
            .I(N__8890));
    InMux I__835 (
            .O(N__8904),
            .I(N__8890));
    InMux I__834 (
            .O(N__8903),
            .I(N__8890));
    InMux I__833 (
            .O(N__8900),
            .I(N__8890));
    InMux I__832 (
            .O(N__8899),
            .I(N__8887));
    LocalMux I__831 (
            .O(N__8890),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__830 (
            .O(N__8887),
            .I(\uu0.l_countZ0Z_1 ));
    InMux I__829 (
            .O(N__8882),
            .I(N__8867));
    InMux I__828 (
            .O(N__8881),
            .I(N__8867));
    InMux I__827 (
            .O(N__8880),
            .I(N__8867));
    InMux I__826 (
            .O(N__8879),
            .I(N__8867));
    InMux I__825 (
            .O(N__8878),
            .I(N__8867));
    LocalMux I__824 (
            .O(N__8867),
            .I(\uu0.l_precountZ0Z_1 ));
    InMux I__823 (
            .O(N__8864),
            .I(N__8854));
    InMux I__822 (
            .O(N__8863),
            .I(N__8854));
    InMux I__821 (
            .O(N__8862),
            .I(N__8854));
    InMux I__820 (
            .O(N__8861),
            .I(N__8851));
    LocalMux I__819 (
            .O(N__8854),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__818 (
            .O(N__8851),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__817 (
            .O(N__8846),
            .I(N__8840));
    InMux I__816 (
            .O(N__8845),
            .I(N__8831));
    InMux I__815 (
            .O(N__8844),
            .I(N__8831));
    InMux I__814 (
            .O(N__8843),
            .I(N__8831));
    InMux I__813 (
            .O(N__8840),
            .I(N__8831));
    LocalMux I__812 (
            .O(N__8831),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__811 (
            .O(N__8828),
            .I(N__8812));
    InMux I__810 (
            .O(N__8827),
            .I(N__8812));
    InMux I__809 (
            .O(N__8826),
            .I(N__8812));
    InMux I__808 (
            .O(N__8825),
            .I(N__8812));
    InMux I__807 (
            .O(N__8824),
            .I(N__8812));
    InMux I__806 (
            .O(N__8823),
            .I(N__8809));
    LocalMux I__805 (
            .O(N__8812),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__804 (
            .O(N__8809),
            .I(\uu0.l_countZ0Z_0 ));
    InMux I__803 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__802 (
            .O(N__8801),
            .I(\uu0.delay_lineZ0Z_1 ));
    InMux I__801 (
            .O(N__8798),
            .I(N__8792));
    InMux I__800 (
            .O(N__8797),
            .I(N__8792));
    LocalMux I__799 (
            .O(N__8792),
            .I(\uu0.delay_lineZ0Z_0 ));
    IoInMux I__798 (
            .O(N__8789),
            .I(N__8786));
    LocalMux I__797 (
            .O(N__8786),
            .I(N__8783));
    Span4Mux_s0_h I__796 (
            .O(N__8783),
            .I(N__8780));
    Odrv4 I__795 (
            .O(N__8780),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__794 (
            .O(N__8777),
            .I(\uu0.un88_ci_3_cascade_ ));
    CascadeMux I__793 (
            .O(N__8774),
            .I(\uu0.un55_ci_cascade_ ));
    InMux I__792 (
            .O(N__8771),
            .I(N__8768));
    LocalMux I__791 (
            .O(N__8768),
            .I(\uu0.un99_ci_0 ));
    CascadeMux I__790 (
            .O(N__8765),
            .I(\uu0.un66_ci_cascade_ ));
    InMux I__789 (
            .O(N__8762),
            .I(N__8747));
    InMux I__788 (
            .O(N__8761),
            .I(N__8747));
    InMux I__787 (
            .O(N__8760),
            .I(N__8747));
    InMux I__786 (
            .O(N__8759),
            .I(N__8747));
    InMux I__785 (
            .O(N__8758),
            .I(N__8747));
    LocalMux I__784 (
            .O(N__8747),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__783 (
            .O(N__8744),
            .I(N__8739));
    CascadeMux I__782 (
            .O(N__8743),
            .I(N__8736));
    InMux I__781 (
            .O(N__8742),
            .I(N__8729));
    InMux I__780 (
            .O(N__8739),
            .I(N__8729));
    InMux I__779 (
            .O(N__8736),
            .I(N__8729));
    LocalMux I__778 (
            .O(N__8729),
            .I(N__8726));
    Odrv4 I__777 (
            .O(N__8726),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    InMux I__776 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__775 (
            .O(N__8720),
            .I(\uu2.un1_l_count_1_2_0 ));
    CascadeMux I__774 (
            .O(N__8717),
            .I(N__8714));
    InMux I__773 (
            .O(N__8714),
            .I(N__8707));
    InMux I__772 (
            .O(N__8713),
            .I(N__8707));
    InMux I__771 (
            .O(N__8712),
            .I(N__8704));
    LocalMux I__770 (
            .O(N__8707),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__769 (
            .O(N__8704),
            .I(\uu2.l_countZ0Z_7 ));
    CascadeMux I__768 (
            .O(N__8699),
            .I(N__8694));
    InMux I__767 (
            .O(N__8698),
            .I(N__8689));
    InMux I__766 (
            .O(N__8697),
            .I(N__8689));
    InMux I__765 (
            .O(N__8694),
            .I(N__8686));
    LocalMux I__764 (
            .O(N__8689),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__763 (
            .O(N__8686),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__762 (
            .O(N__8681),
            .I(N__8678));
    InMux I__761 (
            .O(N__8678),
            .I(N__8673));
    InMux I__760 (
            .O(N__8677),
            .I(N__8668));
    InMux I__759 (
            .O(N__8676),
            .I(N__8668));
    LocalMux I__758 (
            .O(N__8673),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__757 (
            .O(N__8668),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__756 (
            .O(N__8663),
            .I(N__8660));
    InMux I__755 (
            .O(N__8660),
            .I(N__8657));
    LocalMux I__754 (
            .O(N__8657),
            .I(N__8654));
    Odrv4 I__753 (
            .O(N__8654),
            .I(\uu2.un1_l_count_1_3 ));
    CascadeMux I__752 (
            .O(N__8651),
            .I(N__8644));
    InMux I__751 (
            .O(N__8650),
            .I(N__8641));
    InMux I__750 (
            .O(N__8649),
            .I(N__8632));
    InMux I__749 (
            .O(N__8648),
            .I(N__8632));
    InMux I__748 (
            .O(N__8647),
            .I(N__8632));
    InMux I__747 (
            .O(N__8644),
            .I(N__8632));
    LocalMux I__746 (
            .O(N__8641),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__745 (
            .O(N__8632),
            .I(\uu2.l_countZ0Z_2 ));
    CascadeMux I__744 (
            .O(N__8627),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    InMux I__743 (
            .O(N__8624),
            .I(N__8621));
    LocalMux I__742 (
            .O(N__8621),
            .I(\uu2.un1_l_count_2_2 ));
    CascadeMux I__741 (
            .O(N__8618),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    CascadeMux I__740 (
            .O(N__8615),
            .I(\uu2.un350_ci_cascade_ ));
    CascadeMux I__739 (
            .O(N__8612),
            .I(N__8609));
    InMux I__738 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__737 (
            .O(N__8606),
            .I(\uu2.un350_ci ));
    CascadeMux I__736 (
            .O(N__8603),
            .I(N__8598));
    InMux I__735 (
            .O(N__8602),
            .I(N__8591));
    InMux I__734 (
            .O(N__8601),
            .I(N__8591));
    InMux I__733 (
            .O(N__8598),
            .I(N__8591));
    LocalMux I__732 (
            .O(N__8591),
            .I(\uu2.l_countZ0Z_9 ));
    IoInMux I__731 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__730 (
            .O(N__8585),
            .I(N__8582));
    IoSpan4Mux I__729 (
            .O(N__8582),
            .I(N__8579));
    Odrv4 I__728 (
            .O(N__8579),
            .I(clk_in_c));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__22346));
    INV \INVuu2.bitmap_34C  (
            .O(\INVuu2.bitmap_34C_net ),
            .I(N__22357));
    INV \INVuu2.bitmap_218C  (
            .O(\INVuu2.bitmap_218C_net ),
            .I(N__22328));
    INV \INVuu2.bitmap_194C  (
            .O(\INVuu2.bitmap_194C_net ),
            .I(N__22340));
    INV \INVuu2.w_addr_displaying_2_rep1C  (
            .O(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .I(N__22345));
    INV \INVuu2.bitmap_87C  (
            .O(\INVuu2.bitmap_87C_net ),
            .I(N__22351));
    INV \INVuu2.bitmap_203C  (
            .O(\INVuu2.bitmap_203C_net ),
            .I(N__22318));
    INV \INVuu2.w_addr_displaying_fast_7C  (
            .O(\INVuu2.w_addr_displaying_fast_7C_net ),
            .I(N__22327));
    INV \INVuu2.bitmap_90C  (
            .O(\INVuu2.bitmap_90C_net ),
            .I(N__22334));
    INV \INVuu2.w_addr_displaying_fast_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .I(N__22339));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__22309));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__22317));
    INV \INVuu2.bitmap_40C  (
            .O(\INVuu2.bitmap_40C_net ),
            .I(N__22333));
    INV \INVuu2.w_addr_displaying_nesr_8C  (
            .O(\INVuu2.w_addr_displaying_nesr_8C_net ),
            .I(N__22338));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__22344));
    INV \INVuu2.w_addr_user_0C  (
            .O(\INVuu2.w_addr_user_0C_net ),
            .I(N__22350));
    INV \INVuu2.w_addr_user_5C  (
            .O(\INVuu2.w_addr_user_5C_net ),
            .I(N__22356));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__22312));
    INV \INVuu2.w_addr_displaying_4C  (
            .O(\INVuu2.w_addr_displaying_4C_net ),
            .I(N__22337));
    INV \INVuu2.r_data_reg_2C  (
            .O(\INVuu2.r_data_reg_2C_net ),
            .I(N__22335));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__22347));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__10973),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__12176),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__8789),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__14718),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_1_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_1_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_1_6  (
            .in0(N__8959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8992),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_2_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_2_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_1_2_0  (
            .in0(N__8758),
            .in1(N__8986),
            .in2(N__8603),
            .in3(N__9126),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_2_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_2_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_2_1  (
            .in0(N__9013),
            .in1(N__8713),
            .in2(N__8743),
            .in3(N__8760),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_1_2_2 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_1_2_2 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_1_2_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.l_count_8_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8615),
            .in3(N__8697),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22361),
            .ce(),
            .sr(N__22000));
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_2_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_2_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_1_2_3  (
            .in0(N__9127),
            .in1(N__8759),
            .in2(N__8993),
            .in3(N__8601),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_1_2_4 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_1_2_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_1_2_4 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu2.l_count_9_LC_1_2_4  (
            .in0(N__8602),
            .in1(N__8698),
            .in2(N__8612),
            .in3(N__8942),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22361),
            .ce(),
            .sr(N__22000));
    defparam \uu2.l_count_6_LC_1_2_5 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_1_2_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_1_2_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.l_count_6_LC_1_2_5  (
            .in0(N__9014),
            .in1(_gnd_net_),
            .in2(N__8744),
            .in3(N__8761),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22361),
            .ce(),
            .sr(N__22000));
    defparam \uu2.l_count_7_LC_1_2_6 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_1_2_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.l_count_7_LC_1_2_6  (
            .in0(N__8762),
            .in1(N__9015),
            .in2(N__8717),
            .in3(N__8742),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22361),
            .ce(),
            .sr(N__22000));
    defparam \uu2.l_count_3_LC_1_3_0 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_1_3_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_1_3_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uu2.l_count_3_LC_1_3_0  (
            .in0(N__8650),
            .in1(N__8941),
            .in2(N__8681),
            .in3(N__9098),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22359),
            .ce(),
            .sr(N__21997));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_3_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_3_1  (
            .in0(N__8677),
            .in1(N__9154),
            .in2(N__8651),
            .in3(N__9128),
            .lcout(\uu2.un306_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_1_3_2 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_1_3_2 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_1_3_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__9097),
            .in2(_gnd_net_),
            .in3(N__8649),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22359),
            .ce(),
            .sr(N__21997));
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_3_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_3_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_1_3_3  (
            .in0(N__8647),
            .in1(N__8723),
            .in2(N__8663),
            .in3(N__9155),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_3_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_1_3_4  (
            .in0(N__8712),
            .in1(N__8958),
            .in2(N__8699),
            .in3(N__8676),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_1_3_5 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_1_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_1_3_5  (
            .in0(N__8648),
            .in1(N__9156),
            .in2(N__8627),
            .in3(N__8624),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_1_3_6 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_1_3_6 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_1_3_6 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uu2.l_count_4_LC_1_3_6  (
            .in0(_gnd_net_),
            .in1(N__9016),
            .in2(N__8618),
            .in3(N__8990),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22359),
            .ce(),
            .sr(N__21997));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__9295),
            .in2(_gnd_net_),
            .in3(N__9777),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__9439),
            .in2(_gnd_net_),
            .in3(N__9282),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(\uu0.un88_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_9_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_9_3  (
            .in0(N__9491),
            .in1(N__9776),
            .in2(N__8777),
            .in3(N__9418),
            .lcout(\uu0.un110_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_10_1 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_10_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_2_LC_1_10_1  (
            .in0(N__8828),
            .in1(N__8905),
            .in2(_gnd_net_),
            .in3(N__8864),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__9513),
            .sr(N__21990));
    defparam \uu0.l_count_1_LC_1_10_2 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_1_10_2  (
            .in0(N__8904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8827),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__9513),
            .sr(N__21990));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_3  (
            .in0(N__8825),
            .in1(N__8903),
            .in2(_gnd_net_),
            .in3(N__8863),
            .lcout(),
            .ltout(\uu0.un55_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_3_LC_1_10_4 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_10_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \uu0.l_count_3_LC_1_10_4  (
            .in0(N__9570),
            .in1(_gnd_net_),
            .in2(N__8774),
            .in3(N__9401),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__9513),
            .sr(N__21990));
    defparam \uu0.l_count_0_LC_1_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_10_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_10_5  (
            .in0(N__8826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9569),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__9513),
            .sr(N__21990));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_6  (
            .in0(N__8862),
            .in1(N__8824),
            .in2(N__8906),
            .in3(N__9400),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_7_LC_1_10_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_1_10_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_7_LC_1_10_7  (
            .in0(N__8771),
            .in1(N__9419),
            .in2(N__8765),
            .in3(N__9571),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__9513),
            .sr(N__21990));
    defparam \uu0.delay_line_0_LC_1_11_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_11_0  (
            .in0(N__8879),
            .in1(N__9374),
            .in2(N__8924),
            .in3(N__8843),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(N__21992));
    defparam \uu0.l_precount_3_LC_1_11_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_11_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_11_1  (
            .in0(N__8845),
            .in1(N__8922),
            .in2(N__9380),
            .in3(N__8882),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(N__21992));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_11_2 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_11_2  (
            .in0(N__8878),
            .in1(N__9284),
            .in2(N__8923),
            .in3(N__8899),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_1_LC_1_11_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_11_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_precount_1_LC_1_11_3  (
            .in0(N__9375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8880),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(N__21992));
    defparam \uu0.l_precount_2_LC_1_11_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_11_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_1_11_4  (
            .in0(N__8881),
            .in1(N__9376),
            .in2(_gnd_net_),
            .in3(N__8844),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(N__21992));
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_11_5 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI3Q7K1_2_LC_1_11_5  (
            .in0(N__10490),
            .in1(N__8861),
            .in2(N__8846),
            .in3(N__8823),
            .lcout(\uu0.un4_l_count_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_1_LC_1_11_6 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_1_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.delay_line_1_LC_1_11_6  (
            .in0(N__8798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22313),
            .ce(),
            .sr(N__21992));
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_11_7 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_11_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_1_11_7  (
            .in0(N__8804),
            .in1(N__8797),
            .in2(_gnd_net_),
            .in3(N__9556),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_0_LC_1_12_2 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_1_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9363),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22305),
            .ce(),
            .sr(N__21995));
    defparam \buart.Z_rx.hh_0_LC_1_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_13_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9029),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22297),
            .ce(),
            .sr(N__21996));
    defparam \uu2.trig_rd_det_1_LC_2_2_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_2_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_2_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9826),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22360),
            .ce(),
            .sr(N__21973));
    defparam \uu2.l_count_5_LC_2_2_4 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_2_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.l_count_5_LC_2_2_4  (
            .in0(N__9017),
            .in1(N__8960),
            .in2(_gnd_net_),
            .in3(N__8991),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22360),
            .ce(),
            .sr(N__21973));
    defparam \uu2.l_count_0_LC_2_2_7 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_2_2_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_2_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_2_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9132),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22360),
            .ce(),
            .sr(N__21973));
    defparam \uu2.r_addr_5_LC_2_3_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_2_3_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_2_3_0  (
            .in0(N__10133),
            .in1(N__10111),
            .in2(N__10078),
            .in3(N__10211),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \uu2.r_addr_4_LC_2_3_1 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_2_3_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_2_3_1  (
            .in0(N__10110),
            .in1(N__10132),
            .in2(_gnd_net_),
            .in3(N__10210),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \uu2.trig_rd_det_0_LC_2_3_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_2_3_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(N__14870),
            .in2(_gnd_net_),
            .in3(N__10249),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \uu2.vram_rd_clk_LC_2_3_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_2_3_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_2_3_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.vram_rd_clk_LC_2_3_4  (
            .in0(N__14871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8940),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \uu0.sec_clk_LC_2_3_5 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_2_3_5 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_2_3_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(N__14916),
            .in2(_gnd_net_),
            .in3(N__9578),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \uu2.l_count_1_LC_2_3_6 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_2_3_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_2_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_1_LC_2_3_6  (
            .in0(_gnd_net_),
            .in1(N__9158),
            .in2(_gnd_net_),
            .in3(N__9133),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22358),
            .ce(),
            .sr(N__21972));
    defparam \buart.Z_tx.shifter_7_LC_2_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_4_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_4_0  (
            .in0(N__9248),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22352),
            .ce(N__10284),
            .sr(N__21999));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_4_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_4_4  (
            .in0(N__9157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9134),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_0_LC_2_5_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_0_LC_2_5_0  (
            .in0(N__9089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_5_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_1_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9080),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_3_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9071),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_5_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9056),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9050),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_5_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9035),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10409),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_6_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_6_0  (
            .in0(N__9233),
            .in1(N__10596),
            .in2(_gnd_net_),
            .in3(N__9260),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__10595),
            .in2(_gnd_net_),
            .in3(N__9254),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_2_LC_2_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_6_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_6_3  (
            .in0(N__10597),
            .in1(N__9227),
            .in2(_gnd_net_),
            .in3(N__9239),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_3_LC_2_6_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_6_4  (
            .in0(N__9215),
            .in1(N__9164),
            .in2(_gnd_net_),
            .in3(N__10598),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_4_LC_2_6_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_6_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_6_5  (
            .in0(N__10599),
            .in1(N__9203),
            .in2(_gnd_net_),
            .in3(N__9221),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_5_LC_2_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_6_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_6_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_6_6  (
            .in0(N__9182),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(N__9209),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \buart.Z_tx.shifter_6_LC_2_6_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_6_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_6_7  (
            .in0(N__10601),
            .in1(N__9197),
            .in2(_gnd_net_),
            .in3(N__9188),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22342),
            .ce(N__10285),
            .sr(N__21994));
    defparam \uu2.r_data_reg_2_LC_2_7_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_2_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9176),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_2C_net ),
            .ce(N__10405),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_0_LC_2_8_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__9329),
            .in2(_gnd_net_),
            .in3(N__10605),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(N__10286),
            .sr(N__21989));
    defparam \buart.Z_tx.uart_tx_LC_2_8_7 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_8_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_8_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_8_7  (
            .in0(N__10606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9320),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22330),
            .ce(N__10286),
            .sr(N__21989));
    defparam \uu0.l_count_11_LC_2_9_0 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_2_9_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_2_9_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_11_LC_2_9_0  (
            .in0(N__10418),
            .in1(N__9617),
            .in2(N__9809),
            .in3(N__9575),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.l_count_8_LC_2_9_1 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_2_9_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_2_9_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_8_LC_2_9_1  (
            .in0(N__9616),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10484),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.l_count_9_LC_2_9_2 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_2_9_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_2_9_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_9_LC_2_9_2  (
            .in0(N__10485),
            .in1(N__9619),
            .in2(_gnd_net_),
            .in3(N__10449),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.l_count_6_LC_2_9_3 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_2_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_2_9_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_6_LC_2_9_3  (
            .in0(N__9577),
            .in1(N__9494),
            .in2(N__9299),
            .in3(N__9778),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.l_count_5_LC_2_9_4 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_2_9_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_2_9_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_5_LC_2_9_4  (
            .in0(N__9493),
            .in1(N__9440),
            .in2(_gnd_net_),
            .in3(N__9283),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.l_count_13_LC_2_9_6 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_2_9_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_2_9_6 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_13_LC_2_9_6  (
            .in0(N__9848),
            .in1(N__9618),
            .in2(N__9668),
            .in3(N__9576),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22323),
            .ce(N__9512),
            .sr(N__21991));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_10_0 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_10_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_10_0  (
            .in0(N__9878),
            .in1(N__9472),
            .in2(_gnd_net_),
            .in3(N__9649),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_2_10_1 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_2_10_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_15_LC_2_10_1  (
            .in0(N__9621),
            .in1(N__9457),
            .in2(N__9263),
            .in3(N__9560),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__9514),
            .sr(N__21993));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_10_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_10_2  (
            .in0(N__9456),
            .in1(N__9471),
            .in2(N__9885),
            .in3(N__9648),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_10_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_10_3  (
            .in0(N__10444),
            .in1(N__10506),
            .in2(N__9808),
            .in3(N__10479),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_2_10_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_2_10_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_2_10_4  (
            .in0(N__9620),
            .in1(N__9473),
            .in2(N__9497),
            .in3(N__9650),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__9514),
            .sr(N__21993));
    defparam \uu0.l_count_4_LC_2_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_2_10_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_2_10_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu0.l_count_4_LC_2_10_5  (
            .in0(N__9492),
            .in1(N__9438),
            .in2(_gnd_net_),
            .in3(N__9561),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__9514),
            .sr(N__21993));
    defparam \uu0.l_count_10_LC_2_10_6 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_2_10_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_2_10_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu0.l_count_10_LC_2_10_6  (
            .in0(N__10480),
            .in1(N__9622),
            .in2(N__10513),
            .in3(N__10445),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__9514),
            .sr(N__21993));
    defparam \uu0.l_count_RNIGTCU_15_LC_2_10_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNIGTCU_15_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIGTCU_15_LC_2_10_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu0.l_count_RNIGTCU_15_LC_2_10_7  (
            .in0(N__9470),
            .in1(N__10505),
            .in2(N__9458),
            .in3(N__9437),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_11_0  (
            .in0(N__10450),
            .in1(N__9417),
            .in2(N__9701),
            .in3(N__9399),
            .lcout(\uu0.un4_l_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIO2782_16_LC_2_11_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu0.l_count_RNIO2782_16_LC_2_11_1  (
            .in0(N__9386),
            .in1(N__9737),
            .in2(N__9373),
            .in3(N__9640),
            .lcout(),
            .ltout(\uu0.un4_l_count_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_11_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_15_LC_2_11_2  (
            .in0(N__9344),
            .in1(N__9338),
            .in2(N__9332),
            .in3(N__9749),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_11_3 .C_ON=1'b0;
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNIOIDD2_18_LC_2_11_3  (
            .in0(N__9807),
            .in1(N__9679),
            .in2(N__9782),
            .in3(N__9755),
            .lcout(\uu0.un4_l_count_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_2_11_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_2_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_2_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19863),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22306),
            .ce(N__10733),
            .sr(N__21970));
    defparam \resetGen.escKey_5_LC_2_11_5 .C_ON=1'b0;
    defparam \resetGen.escKey_5_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_5_LC_2_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \resetGen.escKey_5_LC_2_11_5  (
            .in0(N__23079),
            .in1(N__22877),
            .in2(N__19878),
            .in3(N__22546),
            .lcout(\resetGen.escKeyZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_2_12_0 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_2_12_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_2_12_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_16_LC_2_12_0  (
            .in0(N__9627),
            .in1(N__9739),
            .in2(N__9722),
            .in3(N__9558),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22298),
            .ce(N__9515),
            .sr(N__21998));
    defparam \uu0.l_count_17_LC_2_12_1 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_12_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_12_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_17_LC_2_12_1  (
            .in0(N__9700),
            .in1(N__9720),
            .in2(N__9743),
            .in3(N__9628),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22298),
            .ce(N__9515),
            .sr(N__21998));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_12_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_12_2  (
            .in0(N__9623),
            .in1(N__9738),
            .in2(N__9721),
            .in3(N__9699),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_12_3 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_12_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_12_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \uu0.l_count_18_LC_2_12_3  (
            .in0(N__9559),
            .in1(_gnd_net_),
            .in2(N__9683),
            .in3(N__9680),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22298),
            .ce(N__9515),
            .sr(N__21998));
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_12_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__9667),
            .in2(_gnd_net_),
            .in3(N__9858),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_12_LC_2_12_6 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_2_12_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_12_LC_2_12_6  (
            .in0(N__9860),
            .in1(N__9887),
            .in2(N__9629),
            .in3(N__9557),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22298),
            .ce(N__9515),
            .sr(N__21998));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_12_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__9886),
            .in2(_gnd_net_),
            .in3(N__9859),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12163),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22291),
            .ce(),
            .sr(N__22001));
    defparam \buart.Z_tx.bitcount_3_LC_4_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_4_2_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_4_2_0 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_4_2_0  (
            .in0(N__11091),
            .in1(N__10570),
            .in2(N__11120),
            .in3(N__10991),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \buart.Z_tx.bitcount_0_LC_4_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_4_2_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_4_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_4_2_1  (
            .in0(N__10569),
            .in1(N__11035),
            .in2(_gnd_net_),
            .in3(N__11090),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \buart.Z_tx.bitcount_2_LC_4_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_4_2_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_4_2_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__10568),
            .in2(_gnd_net_),
            .in3(N__10757),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \uu2.r_addr_2_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_4_2_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_4_2_3  (
            .in0(N__9982),
            .in1(N__10197),
            .in2(N__10015),
            .in3(N__9949),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_4 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(N__9839),
            .in2(_gnd_net_),
            .in3(N__9830),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(\uu2.trig_rd_is_det_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_5 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9812),
            .in3(N__22038),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_1_LC_4_2_6 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_4_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_4_2_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.r_addr_1_LC_4_2_6  (
            .in0(N__9948),
            .in1(_gnd_net_),
            .in2(N__10203),
            .in3(N__9981),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \uu2.r_addr_0_LC_4_2_7 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.r_addr_0_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(N__10193),
            .in2(_gnd_net_),
            .in3(N__9947),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__21981));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_3_0  (
            .in0(_gnd_net_),
            .in1(N__10146),
            .in2(_gnd_net_),
            .in3(N__10040),
            .lcout(),
            .ltout(\uu2.vbuf_raddr.un448_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_3_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_3_1  (
            .in0(N__10171),
            .in1(N__10160),
            .in2(N__10178),
            .in3(N__10125),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__9899),
            .sr(N__21976));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__10076),
            .in2(_gnd_net_),
            .in3(N__10108),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_7_LC_4_3_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_3_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_3_3  (
            .in0(N__10147),
            .in1(N__10041),
            .in2(N__10154),
            .in3(N__10126),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__9899),
            .sr(N__21976));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_3_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_3_4  (
            .in0(N__10007),
            .in1(N__9979),
            .in2(N__9921),
            .in3(N__9945),
            .lcout(\uu2.un404_ci_0 ),
            .ltout(\uu2.un404_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_4_3_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_3_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_3_5  (
            .in0(N__10109),
            .in1(N__10042),
            .in2(N__10082),
            .in3(N__10077),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__9899),
            .sr(N__21976));
    defparam \uu2.r_addr_esr_3_LC_4_3_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_3_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_3_6  (
            .in0(N__10008),
            .in1(N__9980),
            .in2(N__9922),
            .in3(N__9946),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__9899),
            .sr(N__21976));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_4_3_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_4_3_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_4_3_7  (
            .in0(N__14248),
            .in1(N__14387),
            .in2(N__14348),
            .in3(N__14305),
            .lcout(\uu2.un404_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_4_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_4_4_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__10544),
            .in2(_gnd_net_),
            .in3(N__11092),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_4_4_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \uu2.r_data_rdy_LC_4_4_1  (
            .in0(N__22040),
            .in1(N__14882),
            .in2(N__10567),
            .in3(N__10256),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22343),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_2 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_2  (
            .in0(N__15859),
            .in1(N__12352),
            .in2(N__11252),
            .in3(N__15947),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_3 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_3  (
            .in0(N__12353),
            .in1(N__12467),
            .in2(N__15983),
            .in3(N__15860),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_4 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_4  (
            .in0(N__15858),
            .in1(N__15948),
            .in2(N__12566),
            .in3(N__11273),
            .lcout(\uu2.mem0.N_30_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_4_5 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_4_4_5  (
            .in0(N__12482),
            .in1(N__15857),
            .in2(N__15982),
            .in3(N__16787),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_6 .LUT_INIT=16'b1111011010110010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_6  (
            .in0(N__12562),
            .in1(N__11159),
            .in2(N__10220),
            .in3(N__11129),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec2_1_LC_4_5_0 .C_ON=1'b0;
    defparam \Lab_UT.sec2_1_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec2_1_LC_4_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.sec2_1_LC_4_5_0  (
            .in0(N__11813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.sec2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_5_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_5_1 .LUT_INIT=16'b0101010100110000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_4_5_1  (
            .in0(N__12512),
            .in1(N__13497),
            .in2(N__14947),
            .in3(N__11586),
            .lcout(),
            .ltout(\Lab_UT.dispString.m32_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_4_5_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_4_5_2 .LUT_INIT=16'b0001010111111110;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_4_5_2  (
            .in0(N__11481),
            .in1(N__11594),
            .in2(N__10310),
            .in3(N__11326),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_4_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_4_5_3 .LUT_INIT=16'b0001110100110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_4_5_3  (
            .in0(N__10649),
            .in1(N__11584),
            .in2(N__10307),
            .in3(N__11479),
            .lcout(\Lab_UT.dispString.m40_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec1_3_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.sec1_3_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec1_3_LC_4_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec1_3_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11720),
            .lcout(\Lab_UT.sec1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_4_5_5 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_4_5_5  (
            .in0(N__11227),
            .in1(N__11585),
            .in2(N__10298),
            .in3(N__11480),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_4_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_4_5_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__11325),
            .in2(N__10289),
            .in3(N__10331),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min2_0_LC_4_5_7 .C_ON=1'b0;
    defparam \Lab_UT.min2_0_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min2_0_LC_4_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.min2_0_LC_4_5_7  (
            .in0(N__12035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.min2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22336),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_5_LC_4_6_0 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_5_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_5_LC_4_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.alarmchar_5_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12584),
            .lcout(\Lab_UT.alarmcharZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22331),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_4_6_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_4_6_1 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \resetGen.reset_count_4_LC_4_6_1  (
            .in0(N__14675),
            .in1(N__14580),
            .in2(N__10385),
            .in3(N__14548),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22331),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min2_2_LC_4_6_2 .C_ON=1'b0;
    defparam \Lab_UT.min2_2_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min2_2_LC_4_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min2_2_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11984),
            .lcout(\Lab_UT.min2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22331),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_4_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_4_6_3 .LUT_INIT=16'b0101010100110000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_5_LC_4_6_3  (
            .in0(N__10340),
            .in1(N__13498),
            .in2(N__14948),
            .in3(N__11589),
            .lcout(),
            .ltout(\Lab_UT.dispString.m35_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_4_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_4_6_4 .LUT_INIT=16'b0111011101111110;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_4_6_4  (
            .in0(N__11590),
            .in1(N__11327),
            .in2(N__10334),
            .in3(N__11478),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22331),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_4_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_4_6_5 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_4_6_5  (
            .in0(N__11476),
            .in1(N__10316),
            .in2(N__10325),
            .in3(N__11587),
            .lcout(\Lab_UT.dispString.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_4_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_4_6_6 .LUT_INIT=16'b1010001011110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_4_6_6  (
            .in0(N__11588),
            .in1(N__11477),
            .in2(N__14735),
            .in3(N__10373),
            .lcout(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_4_6_7 .C_ON=1'b0;
    defparam \resetGen.rst_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_4_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14579),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22331),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_4_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_4_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dispString.rdy_LC_4_7_0  (
            .in0(N__16336),
            .in1(N__11583),
            .in2(N__11333),
            .in3(N__11475),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec1_2_LC_4_7_1 .C_ON=1'b0;
    defparam \Lab_UT.sec1_2_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec1_2_LC_4_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec1_2_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10672),
            .lcout(\Lab_UT.sec1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec2_0_LC_4_7_2 .C_ON=1'b0;
    defparam \Lab_UT.sec2_0_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec2_0_LC_4_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec2_0_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10751),
            .lcout(\Lab_UT.sec2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_0_LC_4_7_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_0_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_0_LC_4_7_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.alarmchar_0_LC_4_7_3  (
            .in0(N__12755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12878),
            .lcout(\Lab_UT.alarmcharZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_1_LC_4_7_4 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_1_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_1_LC_4_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.alarmchar_1_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__12785),
            .in2(_gnd_net_),
            .in3(N__12754),
            .lcout(\Lab_UT.alarmcharZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_7_5 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_4_7_5  (
            .in0(N__10637),
            .in1(N__11442),
            .in2(N__10367),
            .in3(N__16335),
            .lcout(\Lab_UT.dispString.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min2_1_LC_4_7_6 .C_ON=1'b0;
    defparam \Lab_UT.min2_1_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min2_1_LC_4_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min2_1_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12008),
            .lcout(\Lab_UT.min2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22324),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_4_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_4_7_7 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_4_7_7  (
            .in0(N__10358),
            .in1(N__11441),
            .in2(N__10352),
            .in3(N__11547),
            .lcout(\Lab_UT.dispString.m25_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_0_LC_4_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_4_8_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_4_8_0  (
            .in0(N__11591),
            .in1(N__11473),
            .in2(N__11332),
            .in3(N__16344),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \Lab_UT.didp.regrce2.q_2_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_2_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_2_LC_4_8_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_2_LC_4_8_1  (
            .in0(N__19877),
            .in1(N__20725),
            .in2(N__16391),
            .in3(N__10671),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \Lab_UT.didp.regrce2.q_3_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_3_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_3_LC_4_8_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_3_LC_4_8_2  (
            .in0(N__20726),
            .in1(N__16389),
            .in2(N__19424),
            .in3(N__11716),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \Lab_UT.dictrl.state_0_RNIRNP_1_LC_4_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIRNP_1_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIRNP_1_LC_4_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIRNP_1_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__21453),
            .in2(_gnd_net_),
            .in3(N__21123),
            .lcout(\Lab_UT.dicLdAStens_0 ),
            .ltout(\Lab_UT.dicLdAStens_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_1_LC_4_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_1_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_1_LC_4_8_4 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_1_LC_4_8_4  (
            .in0(N__22768),
            .in1(N__16385),
            .in2(N__10343),
            .in3(N__14752),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \Lab_UT.dispString.cnt_2_LC_4_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_4_8_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_4_8_5  (
            .in0(N__11472),
            .in1(N__11321),
            .in2(_gnd_net_),
            .in3(N__11593),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \Lab_UT.dispString.cnt_1_LC_4_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_4_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_4_8_6  (
            .in0(N__11592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11474),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \buart.Z_tx.bitcount_1_LC_4_8_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_4_8_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_4_8_7 .LUT_INIT=16'b1111100111111100;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_4_8_7  (
            .in0(N__11036),
            .in1(N__11050),
            .in2(N__10607),
            .in3(N__11096),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(),
            .sr(N__21969));
    defparam \buart.Z_rx.bitcount_es_2_LC_4_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_4_9_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_4_9_0 .LUT_INIT=16'b0001010010111110;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_4_9_0  (
            .in0(N__10808),
            .in1(N__10885),
            .in2(N__10859),
            .in3(N__13600),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(N__12119),
            .sr(N__22035));
    defparam \buart.Z_rx.bitcount_es_0_LC_4_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_4_9_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_4_9_1 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_4_9_1  (
            .in0(N__13599),
            .in1(N__10807),
            .in2(N__12648),
            .in3(N__12205),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22307),
            .ce(N__12119),
            .sr(N__22035));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_2  (
            .in0(N__10517),
            .in1(N__10489),
            .in2(_gnd_net_),
            .in3(N__10451),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_9_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_9_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_4_9_3  (
            .in0(N__14831),
            .in1(N__14849),
            .in2(_gnd_net_),
            .in3(N__22034),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_1_LC_4_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_1_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_1_LC_4_9_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m27_1_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__23202),
            .in2(_gnd_net_),
            .in3(N__20414),
            .lcout(\Lab_UT.dictrl.m27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_4_9_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__14519),
            .in2(_gnd_net_),
            .in3(N__14619),
            .lcout(\resetGen.reset_count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_4_10_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_4_10_0  (
            .in0(N__13454),
            .in1(N__10697),
            .in2(N__13340),
            .in3(N__15142),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22299),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.un1_num_5_2_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.un1_num_5_2_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.un1_num_5_2_LC_4_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment3.un1_num_5_2_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__15046),
            .in2(_gnd_net_),
            .in3(N__15229),
            .lcout(),
            .ltout(\Lab_UT.three_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIGRQR1_2_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIGRQR1_2_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIGRQR1_2_LC_4_10_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIGRQR1_2_LC_4_10_2  (
            .in0(N__19874),
            .in1(N__15453),
            .in2(N__10700),
            .in3(N__15141),
            .lcout(\Lab_UT.didp.countrce3.q_5_2 ),
            .ltout(\Lab_UT.didp.countrce3.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_2_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_2_LC_4_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_fast_2_LC_4_10_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_2_LC_4_10_3  (
            .in0(N__10687),
            .in1(N__13453),
            .in2(N__10691),
            .in3(N__13339),
            .lcout(\Lab_UT.didp.countrce3.q_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22299),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_RNII6JA1_2_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_RNII6JA1_2_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_fast_RNII6JA1_2_LC_4_10_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_RNII6JA1_2_LC_4_10_4  (
            .in0(N__11755),
            .in1(N__10750),
            .in2(N__10688),
            .in3(N__11980),
            .lcout(),
            .ltout(\Lab_UT.didp.did_alarmMatch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIQTCC2_2_LC_4_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIQTCC2_2_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIQTCC2_2_LC_4_10_5 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIQTCC2_2_LC_4_10_5  (
            .in0(N__12971),
            .in1(N__10673),
            .in2(N__10652),
            .in3(N__10628),
            .lcout(\Lab_UT.didp.did_alarmMatch_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNISLCD1_1_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNISLCD1_1_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNISLCD1_1_LC_4_10_6 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNISLCD1_1_LC_4_10_6  (
            .in0(N__15230),
            .in1(N__15452),
            .in2(N__15047),
            .in3(N__22766),
            .lcout(\Lab_UT.didp.countrce3.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min2_3_LC_4_10_7 .C_ON=1'b0;
    defparam \Lab_UT.min2_3_LC_4_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min2_3_LC_4_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min2_3_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11944),
            .lcout(\Lab_UT.min2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22299),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min1_1_LC_4_11_0 .C_ON=1'b0;
    defparam \Lab_UT.min1_1_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min1_1_LC_4_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min1_1_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11857),
            .lcout(\Lab_UT.min1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22292),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec2_2_LC_4_11_1 .C_ON=1'b0;
    defparam \Lab_UT.sec2_2_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec2_2_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec2_2_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10627),
            .lcout(\Lab_UT.sec2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22292),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_4_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_4_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__16160),
            .in2(_gnd_net_),
            .in3(N__22037),
            .lcout(\Lab_UT.didp.regrce1.LdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_4_12_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_4_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_0_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16491),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22286),
            .ce(N__10723),
            .sr(N__21974));
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_4_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_4_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_1_LC_4_12_1  (
            .in0(N__22755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22286),
            .ce(N__10723),
            .sr(N__21974));
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_4_12_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_4_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_3_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19419),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22286),
            .ce(N__10723),
            .sr(N__21974));
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_4_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_4_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__10773),
            .in2(_gnd_net_),
            .in3(N__12206),
            .lcout(),
            .ltout(\buart.Z_rx.valid_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_4_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_4_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_4_13_1  (
            .in0(N__10887),
            .in1(N__10841),
            .in2(N__10712),
            .in3(N__10917),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_4_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_4_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_4_13_2  (
            .in0(N__10916),
            .in1(N__10886),
            .in2(N__10844),
            .in3(N__10772),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_1_LC_4_13_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_1_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_1_LC_4_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOUCP_1_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__10837),
            .in2(_gnd_net_),
            .in3(N__10915),
            .lcout(),
            .ltout(\buart.Z_rx.idle_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_4_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_4_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_4_13_4  (
            .in0(N__10888),
            .in1(N__10774),
            .in2(N__10709),
            .in3(N__12207),
            .lcout(\buart.Z_rx.idle ),
            .ltout(\buart.Z_rx.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_1_LC_4_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_1_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_1_LC_4_13_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_1_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10706),
            .in3(N__12136),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(\buart.Z_rx.N_27_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_1_LC_4_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_4_13_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_4_13_6 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_4_13_6  (
            .in0(N__10918),
            .in1(N__10898),
            .in2(N__10703),
            .in3(N__13586),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22281),
            .ce(N__12114),
            .sr(N__22002));
    defparam \buart.Z_rx.bitcount_es_3_LC_4_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_4_13_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_4_13_7 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_4_13_7  (
            .in0(N__13585),
            .in1(N__10797),
            .in2(N__10820),
            .in3(N__10842),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22281),
            .ce(N__12114),
            .sr(N__22002));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_14_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__12208),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_14_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__10919),
            .in2(_gnd_net_),
            .in3(N__10892),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_14_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__10889),
            .in2(_gnd_net_),
            .in3(N__10847),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_14_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__10843),
            .in2(_gnd_net_),
            .in3(N__10811),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_4_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_4_14_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_4_14_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_4_14_4  (
            .in0(N__10798),
            .in1(N__13587),
            .in2(N__10778),
            .in3(N__10781),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22277),
            .ce(N__12115),
            .sr(N__22003));
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23072),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(N__22073),
            .sr(N__22004));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_2_0 .LUT_INIT=16'b1100100111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_5_2_0  (
            .in0(N__11030),
            .in1(N__11002),
            .in2(N__11063),
            .in3(N__11083),
            .lcout(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_2_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_5_2_1  (
            .in0(N__12076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12055),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_2_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__11116),
            .in2(_gnd_net_),
            .in3(N__11029),
            .lcout(\buart.Z_tx.uart_busy_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_2_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_2_4  (
            .in0(N__12054),
            .in1(N__12074),
            .in2(N__12341),
            .in3(N__12257),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(\buart.Z_tx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_2_5 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_2_5  (
            .in0(N__11001),
            .in1(N__11058),
            .in2(N__11105),
            .in3(N__11102),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_2_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_5_2_6  (
            .in0(N__11062),
            .in1(N__11031),
            .in2(N__11006),
            .in3(N__11003),
            .lcout(\buart.Z_tx.un1_bitcount_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_2_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_5_2_7  (
            .in0(N__12075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22349),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_3_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_5_3_1  (
            .in0(N__15979),
            .in1(N__17421),
            .in2(N__14306),
            .in3(N__15837),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_5_3_2 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_5_3_2  (
            .in0(N__15836),
            .in1(N__10969),
            .in2(_gnd_net_),
            .in3(N__15978),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_3_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_5_3_3  (
            .in0(N__15980),
            .in1(N__17492),
            .in2(N__14186),
            .in3(N__15838),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_5_3_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_29_LC_5_3_4  (
            .in0(N__12359),
            .in1(N__12383),
            .in2(_gnd_net_),
            .in3(N__12404),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_3_5 .LUT_INIT=16'b0000001110001001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_19_LC_5_3_5  (
            .in0(N__15977),
            .in1(N__12556),
            .in2(N__11162),
            .in3(N__15835),
            .lcout(\uu2.mem0.w_data_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_6 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_6  (
            .in0(N__15839),
            .in1(N__15981),
            .in2(N__14216),
            .in3(N__17253),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_4_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_36_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__17424),
            .in2(_gnd_net_),
            .in3(N__17486),
            .lcout(\uu2.mem0.bitmap_pmux_sn_N_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_4_1 .LUT_INIT=16'b0100000110111110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_37_LC_5_4_1  (
            .in0(N__17487),
            .in1(N__17912),
            .in2(N__18119),
            .in3(N__17173),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_5_4_2 .LUT_INIT=16'b0001100000000110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_26_LC_5_4_2  (
            .in0(N__17913),
            .in1(N__11141),
            .in2(N__11135),
            .in3(N__18111),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_5_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_5_4_3 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_5_4_3  (
            .in0(N__16969),
            .in1(N__17645),
            .in2(N__11132),
            .in3(N__16127),
            .lcout(\uu2.mem0.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_5_4_4 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_5_4_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_5_4_4  (
            .in0(N__17172),
            .in1(N__18112),
            .in2(N__17921),
            .in3(N__17425),
            .lcout(\uu2.N_34 ),
            .ltout(\uu2.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .LUT_INIT=16'b1010011010100110;
    LogicCell40 \uu2.w_addr_displaying_4_LC_5_4_5  (
            .in0(N__17488),
            .in1(N__17316),
            .in2(N__11123),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__21943));
    defparam \uu2.w_addr_displaying_2_LC_5_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_5_4_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_2_LC_5_4_6  (
            .in0(N__17917),
            .in1(N__17178),
            .in2(N__17321),
            .in3(N__17426),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__21943));
    defparam \uu2.w_addr_displaying_5_LC_5_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_5_4_7 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_5_4_7  (
            .in0(N__17489),
            .in1(N__17320),
            .in2(N__12377),
            .in3(N__17255),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__21943));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_5_5_0 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_5_5_0  (
            .in0(N__11489),
            .in1(N__11168),
            .in2(N__11228),
            .in3(N__11600),
            .lcout(\Lab_UT.dispString.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_4_LC_5_5_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_4_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_4_LC_5_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.un1_w_user_cr_4_LC_5_5_1  (
            .in0(N__11268),
            .in1(N__17073),
            .in2(N__12503),
            .in3(N__11244),
            .lcout(\uu2.un1_w_user_crZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min1_3_LC_5_5_2 .C_ON=1'b0;
    defparam \Lab_UT.min1_3_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min1_3_LC_5_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min1_3_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11831),
            .lcout(\Lab_UT.min1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22332),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_5_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_5_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_5_5_3  (
            .in0(N__15961),
            .in1(N__18113),
            .in2(N__14255),
            .in3(N__15825),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_5_5_4 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_5_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.sec_clkD_LC_5_5_4  (
            .in0(N__14941),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uu0_sec_clkD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22332),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_5_5 .LUT_INIT=16'b0111010101010101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_5_5_5  (
            .in0(N__11192),
            .in1(N__11490),
            .in2(N__11186),
            .in3(N__16346),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_5_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_5_5_6 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__11331),
            .in2(N__11177),
            .in3(N__11174),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22332),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec2_3_LC_5_5_7 .C_ON=1'b0;
    defparam \Lab_UT.sec2_3_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec2_3_LC_5_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec2_3_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11684),
            .lcout(\Lab_UT.sec2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22332),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_6_0 .LUT_INIT=16'b0101100001010000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_5_6_0  (
            .in0(N__11348),
            .in1(N__11639),
            .in2(N__11491),
            .in3(N__16345),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_1 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_5_6_1  (
            .in0(N__11328),
            .in1(_gnd_net_),
            .in2(N__11366),
            .in3(N__11363),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22325),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_6_2 .LUT_INIT=16'b0001110100110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_5_6_2  (
            .in0(N__11354),
            .in1(N__11595),
            .in2(N__11342),
            .in3(N__11482),
            .lcout(\Lab_UT.dispString.m49_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_5_6_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_5_6_3 .LUT_INIT=16'b0000000011010010;
    LogicCell40 \resetGen.reset_count_2_LC_5_6_3  (
            .in0(N__14674),
            .in1(N__14581),
            .in2(N__14621),
            .in3(N__14547),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22325),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_5_6_4  (
            .in0(N__11615),
            .in1(N__11329),
            .in2(_gnd_net_),
            .in3(N__11390),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22325),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec1_0_LC_5_6_5 .C_ON=1'b0;
    defparam \Lab_UT.sec1_0_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec1_0_LC_5_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec1_0_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12716),
            .lcout(\Lab_UT.sec1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22325),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_5_6_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_5_6_6  (
            .in0(N__11606),
            .in1(N__11596),
            .in2(N__11492),
            .in3(N__11330),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22325),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_5_6_7 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_5_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_5_6_7  (
            .in0(N__12463),
            .in1(N__11269),
            .in2(N__12437),
            .in3(N__11245),
            .lcout(\uu2.un1_w_user_lfZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min1_2_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.min1_2_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min1_2_LC_5_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.min1_2_LC_5_7_0  (
            .in0(N__11843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.min1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI8QDI1_2_LC_5_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI8QDI1_2_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI8QDI1_2_LC_5_7_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI8QDI1_2_LC_5_7_1  (
            .in0(N__12711),
            .in1(N__11842),
            .in2(N__20345),
            .in3(N__11751),
            .lcout(\Lab_UT.didp.regrce4.did_alarmMatch_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNIJRBC_1_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNIJRBC_1_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNIJRBC_1_LC_5_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNIJRBC_1_LC_5_7_2  (
            .in0(N__13150),
            .in1(N__13063),
            .in2(_gnd_net_),
            .in3(N__12970),
            .lcout(\Lab_UT.didp.countrce2.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_2_LC_5_7_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_2_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_2_LC_5_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.alarmchar_2_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12599),
            .lcout(\Lab_UT.alarmcharZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.min1_0_LC_5_7_4 .C_ON=1'b0;
    defparam \Lab_UT.min1_0_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.min1_0_LC_5_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.min1_0_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11876),
            .lcout(\Lab_UT.min1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_5 .LUT_INIT=16'b0110010001000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_5  (
            .in0(N__11633),
            .in1(N__11471),
            .in2(N__11624),
            .in3(N__16337),
            .lcout(\Lab_UT.dispString.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_6_LC_5_7_6 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_6_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_6_LC_5_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.alarmchar_6_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12722),
            .lcout(\Lab_UT.alarmcharZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22316),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_7_7 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_5_7_7  (
            .in0(N__11582),
            .in1(N__11513),
            .in2(N__11507),
            .in3(N__11470),
            .lcout(\Lab_UT.dispString.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_5_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_5_8_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_5_8_0  (
            .in0(N__15223),
            .in1(N__11875),
            .in2(N__20140),
            .in3(N__12031),
            .lcout(),
            .ltout(\Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRSKRA_0_LC_5_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRSKRA_0_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRSKRA_0_LC_5_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIRSKRA_0_LC_5_8_1  (
            .in0(N__11384),
            .in1(N__11378),
            .in2(N__11369),
            .in3(N__11645),
            .lcout(\Lab_UT.alarmMatch ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_fast_0_LC_5_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_fast_0_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_fast_0_LC_5_8_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce2.q_fast_0_LC_5_8_2  (
            .in0(N__13277),
            .in1(N__12092),
            .in2(N__11759),
            .in3(N__13791),
            .lcout(\Lab_UT.didp.q_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNIUST81_3_LC_5_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNIUST81_3_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNIUST81_3_LC_5_8_3 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNIUST81_3_LC_5_8_3  (
            .in0(N__11732),
            .in1(N__19423),
            .in2(N__18716),
            .in3(N__13004),
            .lcout(\Lab_UT.didp.countrce2.q_5_3 ),
            .ltout(\Lab_UT.didp.countrce2.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_fast_3_LC_5_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_fast_3_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_fast_3_LC_5_8_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.didp.countrce2.q_fast_3_LC_5_8_4  (
            .in0(N__13278),
            .in1(N__11699),
            .in2(N__11723),
            .in3(N__13792),
            .lcout(\Lab_UT.didp.countrce2.q_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_fast_RNIOS8A1_3_LC_5_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_fast_RNIOS8A1_3_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_fast_RNIOS8A1_3_LC_5_8_5 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \Lab_UT.didp.countrce2.q_fast_RNIOS8A1_3_LC_5_8_5  (
            .in0(N__11715),
            .in1(N__11695),
            .in2(_gnd_net_),
            .in3(N__11683),
            .lcout(\Lab_UT.didp.did_alarmMatch_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_5_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_5_8_6 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_5_8_6  (
            .in0(N__13005),
            .in1(N__13790),
            .in2(N__13283),
            .in3(N__11660),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_5_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_5_8_7 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_5_8_7  (
            .in0(N__12091),
            .in1(N__13279),
            .in2(N__13793),
            .in3(N__13068),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22308),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_9_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_9_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_RNINLQC1_1_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_RNINLQC1_1_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_fast_RNINLQC1_1_LC_5_9_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_RNINLQC1_1_LC_5_9_1  (
            .in0(N__11773),
            .in1(N__11858),
            .in2(N__12904),
            .in3(N__12004),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_RNI077E5_1_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_RNI077E5_1_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_fast_RNI077E5_1_LC_5_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_RNI077E5_1_LC_5_9_2  (
            .in0(N__11654),
            .in1(N__11795),
            .in2(N__11648),
            .in3(N__11882),
            .lcout(\Lab_UT.didp.did_alarmMatch_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.un1_num_5_2_LC_5_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment2.un1_num_5_2_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__13133),
            .in2(_gnd_net_),
            .in3(N__13064),
            .lcout(),
            .ltout(\Lab_UT.three_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_5_9_4 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_5_9_4  (
            .in0(N__18704),
            .in1(N__19872),
            .in2(N__11816),
            .in3(N__12959),
            .lcout(\Lab_UT.didp.countrce2.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_fast_RNIIM8A1_1_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_fast_RNIIM8A1_1_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_fast_RNIIM8A1_1_LC_5_9_5 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \Lab_UT.didp.countrce2.q_fast_RNIIM8A1_1_LC_5_9_5  (
            .in0(N__11785),
            .in1(N__14751),
            .in2(_gnd_net_),
            .in3(N__11812),
            .lcout(\Lab_UT.didp.did_alarmMatch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_fast_1_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_fast_1_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_fast_1_LC_5_9_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce2.q_fast_1_LC_5_9_6  (
            .in0(N__13274),
            .in1(N__12695),
            .in2(N__11789),
            .in3(N__13776),
            .lcout(\Lab_UT.didp.countrce2.q_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22300),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_5_9_7 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_5_9_7  (
            .in0(N__12694),
            .in1(N__13275),
            .in2(N__13786),
            .in3(N__13134),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22300),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_1_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_1_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_fast_1_LC_5_10_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_1_LC_5_10_0  (
            .in0(N__13449),
            .in1(N__13327),
            .in2(N__13181),
            .in3(N__11774),
            .lcout(\Lab_UT.didp.countrce3.q_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22293),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_fast_3_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_fast_3_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_fast_3_LC_5_10_1 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \Lab_UT.didp.countrce4.q_fast_3_LC_5_10_1  (
            .in0(N__11893),
            .in1(N__13396),
            .in2(N__13226),
            .in3(N__13192),
            .lcout(\Lab_UT.didp.q_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22293),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIMAAB1_2_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIMAAB1_2_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIMAAB1_2_LC_5_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIMAAB1_2_LC_5_10_2  (
            .in0(N__15139),
            .in1(N__15033),
            .in2(_gnd_net_),
            .in3(N__15219),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNI529A2_3_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNI529A2_3_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNI529A2_3_LC_5_10_3 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNI529A2_3_LC_5_10_3  (
            .in0(N__15086),
            .in1(N__19414),
            .in2(N__11762),
            .in3(N__15454),
            .lcout(\Lab_UT.didp.countrce3.q_5_3 ),
            .ltout(\Lab_UT.didp.countrce3.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_3_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_3_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_fast_3_LC_5_10_4 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_3_LC_5_10_4  (
            .in0(N__13450),
            .in1(N__13328),
            .in2(N__11906),
            .in3(N__11903),
            .lcout(\Lab_UT.didp.countrce3.q_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22293),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_fast_RNIVTQC1_3_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_fast_RNIVTQC1_3_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_fast_RNIVTQC1_3_LC_5_10_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.countrce3.q_fast_RNIVTQC1_3_LC_5_10_5  (
            .in0(N__11902),
            .in1(N__11827),
            .in2(N__11894),
            .in3(N__11943),
            .lcout(\Lab_UT.didp.countrce3.did_alarmMatch_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_5_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_5_10_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_5_10_6  (
            .in0(N__13397),
            .in1(N__13508),
            .in2(N__20123),
            .in3(N__13221),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22293),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.un1_num_11_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.un1_num_11_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.un1_num_11_LC_5_10_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.bcd2segment3.un1_num_11_LC_5_10_7  (
            .in0(N__15220),
            .in1(N__15140),
            .in2(N__15109),
            .in3(N__15032),
            .lcout(\Lab_UT.nine_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_5_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_0_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16489),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22287),
            .ce(N__13478),
            .sr(N__21975));
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_5_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_1_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22767),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22287),
            .ce(N__13478),
            .sr(N__21975));
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_5_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_2_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19876),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22287),
            .ce(N__13478),
            .sr(N__21975));
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_5_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_3_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19407),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22287),
            .ce(N__13478),
            .sr(N__21975));
    defparam \Lab_UT.didp.ce_11_2_LC_5_12_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_11_2_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_11_2_LC_5_12_0 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \Lab_UT.didp.ce_11_2_LC_5_12_0  (
            .in0(N__15440),
            .in1(N__21429),
            .in2(N__15377),
            .in3(N__20655),
            .lcout(\Lab_UT.didp.ce_11_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_RNI0RGF_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNI0RGF_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNI0RGF_LC_5_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNI0RGF_LC_5_12_1  (
            .in0(N__21430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15376),
            .lcout(\Lab_UT.dicLdAMones_0 ),
            .ltout(\Lab_UT.dicLdAMones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_0_LC_5_12_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_0_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_0_LC_5_12_2 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \Lab_UT.didp.regrce3.q_0_LC_5_12_2  (
            .in0(N__16493),
            .in1(N__20657),
            .in2(N__12038),
            .in3(N__12027),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(),
            .sr(N__21977));
    defparam \Lab_UT.didp.regrce3.q_1_LC_5_12_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_1_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_1_LC_5_12_3 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_1_LC_5_12_3  (
            .in0(N__22706),
            .in1(N__11955),
            .in2(N__20666),
            .in3(N__12003),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(),
            .sr(N__21977));
    defparam \Lab_UT.didp.regrce3.q_2_LC_5_12_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_2_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_2_LC_5_12_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \Lab_UT.didp.regrce3.q_2_LC_5_12_4  (
            .in0(N__19875),
            .in1(N__20658),
            .in2(N__11960),
            .in3(N__11979),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(),
            .sr(N__21977));
    defparam \Lab_UT.didp.regrce3.q_3_LC_5_12_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_3_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_3_LC_5_12_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_3_LC_5_12_5  (
            .in0(N__20656),
            .in1(N__19402),
            .in2(N__11945),
            .in3(N__11959),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(),
            .sr(N__21977));
    defparam \resetGen.escKey_4_LC_5_12_6 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_5_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \resetGen.escKey_4_LC_5_12_6  (
            .in0(N__16492),
            .in1(N__22705),
            .in2(N__19418),
            .in3(N__22460),
            .lcout(),
            .ltout(\resetGen.escKeyZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_5_12_7 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_5_12_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \resetGen.escKey_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__11921),
            .in2(N__11909),
            .in3(N__12135),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_13_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_5_13_0  (
            .in0(N__13580),
            .in1(N__13637),
            .in2(N__13627),
            .in3(N__13651),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_13_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_5_13_1  (
            .in0(N__13723),
            .in1(N__13581),
            .in2(_gnd_net_),
            .in3(N__13738),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_13_2 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_5_13_2  (
            .in0(N__13690),
            .in1(N__13628),
            .in2(N__13598),
            .in3(N__13676),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22278),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_5_13_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_5_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_5_13_3  (
            .in0(N__13666),
            .in1(N__13689),
            .in2(N__13528),
            .in3(N__13737),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_5_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_5_13_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__13650),
            .in2(N__12224),
            .in3(N__13722),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_13_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__12221),
            .in2(N__12215),
            .in3(N__12212),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_13_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_5_13_6  (
            .in0(N__13867),
            .in1(N__12164),
            .in2(_gnd_net_),
            .in3(N__12148),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(\buart.Z_rx.startbit_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_13_7 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_5_13_7  (
            .in0(N__12149),
            .in1(N__13619),
            .in2(N__12140),
            .in3(N__12137),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI5RHS_0_LC_5_14_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI5RHS_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI5RHS_0_LC_5_14_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI5RHS_0_LC_5_14_7  (
            .in0(N__18712),
            .in1(N__16450),
            .in2(_gnd_net_),
            .in3(N__13084),
            .lcout(\Lab_UT.didp.countrce2.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIINVH_2_LC_6_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_6_1_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu2.w_addr_user_RNIINVH_2_LC_6_1_6  (
            .in0(N__14332),
            .in1(N__13907),
            .in2(N__14177),
            .in3(N__12302),
            .lcout(\uu2.un3_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_2_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__12077),
            .in2(N__12059),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_2_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__12266),
            .in2(_gnd_net_),
            .in3(N__12041),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__22341),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_2_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_6_2_2  (
            .in0(N__12315),
            .in1(N__12340),
            .in2(_gnd_net_),
            .in3(N__12326),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__22341),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_2_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__12287),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__22341),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_2_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_6_2_4  (
            .in0(N__12316),
            .in1(N__12296),
            .in2(_gnd_net_),
            .in3(N__12320),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__22341),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_2_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_6_2_5  (
            .in0(N__12277),
            .in1(N__12317),
            .in2(_gnd_net_),
            .in3(N__12305),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22341),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_6_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_6_2_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.w_addr_user_nesr_RNI9006_8_LC_6_2_6  (
            .in0(N__14085),
            .in1(N__14483),
            .in2(_gnd_net_),
            .in3(N__14283),
            .lcout(\uu2.un3_w_addr_user_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_2_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_2_7  (
            .in0(N__12295),
            .in1(N__12286),
            .in2(N__12278),
            .in3(N__12265),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_6_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_6_3_0 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_6_3_0  (
            .in0(N__16118),
            .in1(N__14086),
            .in2(N__15856),
            .in3(N__15988),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_3_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_3_1 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_6_3_1  (
            .in0(N__17920),
            .in1(N__14370),
            .in2(N__15995),
            .in3(N__15844),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_6_3_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_6_3_2 .LUT_INIT=16'b1000000100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_44_LC_6_3_2  (
            .in0(N__17558),
            .in1(N__17919),
            .in2(N__18118),
            .in3(N__13988),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3  (
            .in0(N__15987),
            .in1(N__17174),
            .in2(N__14341),
            .in3(N__15840),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_6_3_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_6_3_5 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_31_LC_6_3_5  (
            .in0(N__17249),
            .in1(N__16970),
            .in2(N__15689),
            .in3(N__16117),
            .lcout(\uu2.mem0.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_51_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__17476),
            .in2(_gnd_net_),
            .in3(N__17765),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_6_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_6_3_7 .LUT_INIT=16'b1010001010101000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_43_LC_6_3_7  (
            .in0(N__16801),
            .in1(N__18104),
            .in2(N__12386),
            .in3(N__17557),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_6_4_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.rdy_RNIGIDK3_LC_6_4_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dispString.rdy_RNIGIDK3_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__15984),
            .in2(_gnd_net_),
            .in3(N__15803),
            .lcout(N_272_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI17I72_5_LC_6_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI17I72_5_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI17I72_5_LC_6_4_2 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \uu2.w_addr_displaying_RNI17I72_5_LC_6_4_2  (
            .in0(N__17491),
            .in1(_gnd_net_),
            .in2(N__12376),
            .in3(N__17254),
            .lcout(\uu2.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_4_3 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_42_LC_6_4_3  (
            .in0(N__17171),
            .in1(N__17422),
            .in2(_gnd_net_),
            .in3(N__17490),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIB2283_5_LC_6_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIB2283_5_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIB2283_5_LC_6_4_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIB2283_5_LC_6_4_4  (
            .in0(N__15741),
            .in1(N__12526),
            .in2(_gnd_net_),
            .in3(N__18296),
            .lcout(\uu2.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIEHP31_6_LC_6_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIEHP31_6_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIEHP31_6_LC_6_4_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIEHP31_6_LC_6_4_6  (
            .in0(N__15681),
            .in1(N__16968),
            .in2(_gnd_net_),
            .in3(N__16121),
            .lcout(\uu2.N_57 ),
            .ltout(\uu2.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_1_LC_6_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_1_LC_6_4_7 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIFOBB3_1_LC_6_4_7  (
            .in0(N__12525),
            .in1(N__17918),
            .in2(N__12569),
            .in3(N__17423),
            .lcout(\uu2.w_data_i_a3_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_5_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_21_LC_6_5_0  (
            .in0(N__17396),
            .in1(_gnd_net_),
            .in2(N__15748),
            .in3(N__12527),
            .lcout(),
            .ltout(\uu2.mem0.w_data_0_a3_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_1  (
            .in0(N__15993),
            .in1(N__12502),
            .in2(N__12545),
            .in3(N__15828),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNITJLE1_5_LC_6_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNITJLE1_5_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNITJLE1_5_LC_6_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNITJLE1_5_LC_6_5_2  (
            .in0(N__17485),
            .in1(N__17180),
            .in2(N__18116),
            .in3(N__17248),
            .lcout(\uu2.w_data_displaying_2_i_a2_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_4_LC_6_5_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_4_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_4_LC_6_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.alarmchar_4_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12593),
            .lcout(\Lab_UT.alarmcharZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22320),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_0_LC_6_5_4 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_0_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_0_LC_6_5_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.un1_w_user_lf_0_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__12480),
            .in2(_gnd_net_),
            .in3(N__12501),
            .lcout(\uu2.un1_w_user_lf_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_LC_6_5_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_LC_6_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.un1_w_user_cr_LC_6_5_5  (
            .in0(N__12481),
            .in1(N__12462),
            .in2(N__12436),
            .in3(N__12446),
            .lcout(uu2_un1_w_user_cr_0),
            .ltout(uu2_un1_w_user_cr_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_5_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_5_6 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__15992),
            .in2(N__12440),
            .in3(N__12432),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIGEPH1_2_LC_6_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIGEPH1_2_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIGEPH1_2_LC_6_5_7 .LUT_INIT=16'b0110101000001000;
    LogicCell40 \uu2.w_addr_displaying_RNIGEPH1_2_LC_6_5_7  (
            .in0(N__17179),
            .in1(N__17395),
            .in2(N__18103),
            .in3(N__17484),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_2_LC_6_6_0 .LUT_INIT=16'b0111011011110111;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_2_LC_6_6_0  (
            .in0(N__12968),
            .in1(N__13017),
            .in2(N__13102),
            .in3(N__13156),
            .lcout(\Lab_UT.bcd2segment2.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_4_LC_6_6_1 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_4_LC_6_6_1  (
            .in0(N__13151),
            .in1(N__13085),
            .in2(N__13022),
            .in3(N__12963),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_5_LC_6_6_2 .LUT_INIT=16'b1111110110011000;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_5_LC_6_6_2  (
            .in0(N__12964),
            .in1(N__13009),
            .in2(N__13100),
            .in3(N__13152),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_6_LC_6_6_3 .LUT_INIT=16'b1111100010100101;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_6_LC_6_6_3  (
            .in0(N__13153),
            .in1(N__13089),
            .in2(N__13023),
            .in3(N__12965),
            .lcout(\Lab_UT.bcd2segment2.segmentUQ_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_6_6_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_0_LC_6_6_4 .LUT_INIT=16'b1011111101101101;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_0_LC_6_6_4  (
            .in0(N__12966),
            .in1(N__13013),
            .in2(N__13101),
            .in3(N__13154),
            .lcout(\Lab_UT.bcd2segment2.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_6_6_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_0_1_LC_6_6_5 .LUT_INIT=16'b0100100101111111;
    LogicCell40 \Lab_UT.bcd2segment2.segment_0_1_LC_6_6_5  (
            .in0(N__13155),
            .in1(N__13093),
            .in2(N__13024),
            .in3(N__12967),
            .lcout(\Lab_UT.bcd2segment2.segment_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_6_6_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_3_LC_6_6_6 .LUT_INIT=16'b1110110011011010;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_3_LC_6_6_6  (
            .in0(N__12969),
            .in1(N__13018),
            .in2(N__13103),
            .in3(N__13157),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_6_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_6_6_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_308_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12572),
            .in3(N__20058),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__21940));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_64_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_64_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__G_64_LC_6_7_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__G_64_LC_6_7_0  (
            .in0(N__12850),
            .in1(N__12803),
            .in2(N__14790),
            .in3(N__14722),
            .lcout(\Lab_UT.dictrl.G_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_6_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_0_LC_6_7_1  (
            .in0(N__12657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22304),
            .ce(N__12623),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m6_xx_mm_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m6_xx_mm_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m6_xx_mm_LC_6_7_2 .LUT_INIT=16'b0000000011001110;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__m6_xx_mm_LC_6_7_2  (
            .in0(N__12614),
            .in1(N__12743),
            .in2(N__12781),
            .in3(N__16415),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_7_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_7_3  (
            .in0(N__12742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12773),
            .lcout(),
            .ltout(\Lab_UT.dictrl.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_7_4 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_7_4  (
            .in0(N__12613),
            .in1(N__12867),
            .in2(N__12605),
            .in3(N__16414),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1_0 ),
            .ltout(\Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNINRI3E_0_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNINRI3E_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNINRI3E_0_LC_6_7_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNINRI3E_0_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__14774),
            .in2(N__12602),
            .in3(N__12823),
            .lcout(\Lab_UT.dictrl.next_alarmstate_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNIT8JUD_0_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIT8JUD_0_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIT8JUD_0_LC_6_7_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNIT8JUD_0_LC_6_7_6  (
            .in0(N__14775),
            .in1(_gnd_net_),
            .in2(N__12830),
            .in3(N__12802),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_7_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_7_7  (
            .in0(N__12744),
            .in1(_gnd_net_),
            .in2(N__12874),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmchar9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_6_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_6_8_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_1_LC_6_8_0  (
            .in0(N__14794),
            .in1(N__12852),
            .in2(_gnd_net_),
            .in3(N__12805),
            .lcout(\Lab_UT.alarmchar10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_6_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_6_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_6_8_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_2_LC_6_8_1  (
            .in0(N__12806),
            .in1(N__14795),
            .in2(_gnd_net_),
            .in3(N__12853),
            .lcout(\Lab_UT.alarmchar10_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_6_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_6_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_0_LC_6_8_2  (
            .in0(N__14791),
            .in1(N__12827),
            .in2(_gnd_net_),
            .in3(N__12851),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_6_8_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_6_8_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_LC_6_8_3  (
            .in0(N__12829),
            .in1(N__14793),
            .in2(_gnd_net_),
            .in3(N__12854),
            .lcout(\Lab_UT.dictrl.alarmstate_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_6_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_6_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_1_LC_6_8_4  (
            .in0(N__14792),
            .in1(N__12828),
            .in2(_gnd_net_),
            .in3(N__12804),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_6_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_6_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__12777),
            .in2(_gnd_net_),
            .in3(N__12745),
            .lcout(\Lab_UT.alarmchar_2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_8_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_8_6  (
            .in0(N__15455),
            .in1(N__16474),
            .in2(_gnd_net_),
            .in3(N__15221),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_0_LC_6_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_0_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_0_LC_6_8_7 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_0_LC_6_8_7  (
            .in0(N__16475),
            .in1(N__20727),
            .in2(N__16390),
            .in3(N__12712),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22295),
            .ce(),
            .sr(N__21971));
    defparam \Lab_UT.didp.countrce2.q_RNINQL01_1_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNINQL01_1_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNINQL01_1_LC_6_9_0 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNINQL01_1_LC_6_9_0  (
            .in0(N__13062),
            .in1(N__13132),
            .in2(N__18705),
            .in3(N__22737),
            .lcout(\Lab_UT.didp.countrce2.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_6_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment1.un1_num_5_2_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__18344),
            .in2(_gnd_net_),
            .in3(N__18462),
            .lcout(\Lab_UT.three_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_6_9_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_6_9_2  (
            .in0(N__12958),
            .in1(N__13764),
            .in2(N__12686),
            .in3(N__13276),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22289),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_9_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_6_9_3  (
            .in0(N__13451),
            .in1(N__12677),
            .in2(N__13335),
            .in3(N__15222),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22289),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_6_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.bcd2segment1.un1_num_11_LC_6_9_4  (
            .in0(N__18523),
            .in1(N__18481),
            .in2(N__18364),
            .in3(N__18395),
            .lcout(\Lab_UT.nine ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_9_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__13713),
            .in2(_gnd_net_),
            .in3(N__13601),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22289),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_6_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_6_9_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_6_9_6  (
            .in0(N__13326),
            .in1(N__13180),
            .in2(N__15042),
            .in3(N__13452),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22289),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.un1_num_7_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.un1_num_7_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.un1_num_7_LC_6_9_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.bcd2segment2.un1_num_7_LC_6_9_7  (
            .in0(N__13131),
            .in1(N__13061),
            .in2(N__13025),
            .in3(N__12957),
            .lcout(\Lab_UT.five ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_6_10_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_6_10_0  (
            .in0(N__13448),
            .in1(N__12911),
            .in2(N__13334),
            .in3(N__15087),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_fast_1_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_fast_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_fast_1_LC_6_10_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_fast_1_LC_6_10_1  (
            .in0(N__13387),
            .in1(N__12887),
            .in2(N__12905),
            .in3(N__13220),
            .lcout(\Lab_UT.didp.q_fast_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNI33OG1_1_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNI33OG1_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNI33OG1_1_LC_6_10_2 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNI33OG1_1_LC_6_10_2  (
            .in0(N__20110),
            .in1(N__18938),
            .in2(N__20184),
            .in3(N__22736),
            .lcout(\Lab_UT.didp.countrce4.q_5_1 ),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_6_10_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_6_10_3  (
            .in0(N__13388),
            .in1(N__13215),
            .in2(N__12881),
            .in3(N__20178),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_10_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_6_10_4  (
            .in0(N__13193),
            .in1(N__13390),
            .in2(N__13225),
            .in3(N__20242),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.un1_num_5_2_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.un1_num_5_2_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.un1_num_5_2_LC_6_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment4.un1_num_5_2_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__20177),
            .in2(_gnd_net_),
            .in3(N__20111),
            .lcout(),
            .ltout(\Lab_UT.three_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_10_6 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_10_6  (
            .in0(N__19856),
            .in1(N__18939),
            .in2(N__13238),
            .in3(N__20316),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_10_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_6_10_7  (
            .in0(N__13389),
            .in1(N__20312),
            .in2(N__13235),
            .in3(N__13216),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22285),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_1_3_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_1_3_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_1_3_LC_6_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.reset_RNO_1_3_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__20240),
            .in2(_gnd_net_),
            .in3(N__20173),
            .lcout(),
            .ltout(\Lab_UT.didp.reset_12_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_6_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_6_11_1  (
            .in0(N__16292),
            .in1(N__20109),
            .in2(N__13232),
            .in3(N__20311),
            .lcout(),
            .ltout(\Lab_UT.didp.reset_12_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_6_11_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_6_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_6_11_2  (
            .in0(N__13847),
            .in1(N__13359),
            .in2(N__13229),
            .in3(N__13817),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(),
            .sr(N__21978));
    defparam \Lab_UT.didp.countrce4.q_RNIPP8Q_1_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNIPP8Q_1_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNIPP8Q_1_LC_6_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNIPP8Q_1_LC_6_11_3  (
            .in0(N__20172),
            .in1(N__20107),
            .in2(_gnd_net_),
            .in3(N__20310),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNIEP822_3_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNIEP822_3_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNIEP822_3_LC_6_11_4 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNIEP822_3_LC_6_11_4  (
            .in0(N__18934),
            .in1(N__19406),
            .in2(N__13196),
            .in3(N__20241),
            .lcout(\Lab_UT.didp.countrce4.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_0_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_6_11_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_6_11_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_6_11_5  (
            .in0(N__16293),
            .in1(N__13846),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(),
            .sr(N__21978));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_11_6 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_11_6  (
            .in0(N__20108),
            .in1(_gnd_net_),
            .in2(N__18941),
            .in3(N__16488),
            .lcout(\Lab_UT.didp.countrce4.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_6_11_7 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_6_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__13502),
            .in2(_gnd_net_),
            .in3(N__14945),
            .lcout(oneSecStrb),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_6_12_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_6_12_0  (
            .in0(N__21127),
            .in1(N__15352),
            .in2(N__20665),
            .in3(N__22039),
            .lcout(\Lab_UT.didp.regrce4.LdAMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.un26_ce_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.un26_ce_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.un26_ce_LC_6_12_1 .LUT_INIT=16'b0100110000001100;
    LogicCell40 \Lab_UT.didp.un26_ce_LC_6_12_1  (
            .in0(N__13842),
            .in1(N__13465),
            .in2(N__13820),
            .in3(N__18646),
            .lcout(\Lab_UT.didp.un26_ce_0 ),
            .ltout(\Lab_UT.didp.un26_ce_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_2_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_6_12_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \Lab_UT.didp.ce_2_LC_6_12_2  (
            .in0(N__13466),
            .in1(_gnd_net_),
            .in2(N__13457),
            .in3(N__16316),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(N__21982));
    defparam \Lab_UT.didp.ce_RNO_0_3_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNO_0_3_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNO_0_3_LC_6_12_3 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \Lab_UT.didp.ce_RNO_0_3_LC_6_12_3  (
            .in0(N__18940),
            .in1(N__20654),
            .in2(N__15353),
            .in3(N__21128),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_3_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_6_12_4 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \Lab_UT.didp.ce_3_LC_6_12_4  (
            .in0(N__16299),
            .in1(N__13360),
            .in2(N__13406),
            .in3(N__13403),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(N__21982));
    defparam \Lab_UT.didp.reset_2_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_6_12_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_6_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_6_12_5  (
            .in0(N__13845),
            .in1(N__13819),
            .in2(N__13364),
            .in3(N__16301),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(N__21982));
    defparam \Lab_UT.didp.ce_1_LC_6_12_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_6_12_6 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \Lab_UT.didp.ce_1_LC_6_12_6  (
            .in0(N__18647),
            .in1(N__16317),
            .in2(_gnd_net_),
            .in3(N__13843),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(N__21982));
    defparam \Lab_UT.didp.reset_1_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_6_12_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_6_12_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_6_12_7  (
            .in0(N__13844),
            .in1(N__13818),
            .in2(_gnd_net_),
            .in3(N__16300),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22276),
            .ce(),
            .sr(N__21982));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_13_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__13739),
            .in2(N__13724),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_13_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__13691),
            .in2(_gnd_net_),
            .in3(N__13670),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_13_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_6_13_2  (
            .in0(N__13589),
            .in1(N__13667),
            .in2(_gnd_net_),
            .in3(N__13655),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__22272),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_13_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__13652),
            .in2(_gnd_net_),
            .in3(N__13631),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_13_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_6_13_4  (
            .in0(N__13623),
            .in1(N__13588),
            .in2(N__13529),
            .in3(N__13532),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22272),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_19_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_19_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_19_LC_6_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_19_LC_6_13_5  (
            .in0(N__21126),
            .in1(N__15470),
            .in2(_gnd_net_),
            .in3(N__13853),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_2_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_2_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_2_LC_6_13_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_2_LC_6_13_6  (
            .in0(N__21452),
            .in1(N__20663),
            .in2(N__13511),
            .in3(N__15497),
            .lcout(\Lab_UT.dictrl.N_11_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_3_LC_6_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_3_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_3_LC_6_14_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_1_3_LC_6_14_0  (
            .in0(N__13898),
            .in1(N__15518),
            .in2(N__13886),
            .in3(N__15487),
            .lcout(\Lab_UT.dictrl.g0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_LC_6_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_6_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_6_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13875),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22270),
            .ce(N__22071),
            .sr(N__22005));
    defparam \buart.Z_rx.shifter_fast_7_LC_6_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_6_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_6_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_6_14_5  (
            .in0(N__13877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22270),
            .ce(N__22071),
            .sr(N__22005));
    defparam \buart.Z_rx.shifter_7_rep1_LC_6_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_6_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13876),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22270),
            .ce(N__22071),
            .sr(N__22005));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_22_LC_6_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_22_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_22_LC_6_14_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_22_LC_6_14_7  (
            .in0(N__23033),
            .in1(N__22876),
            .in2(N__16874),
            .in3(N__22558),
            .lcout(\Lab_UT.dictrl.g2_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_6_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_6_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_6_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22727),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__22069),
            .sr(N__22006));
    defparam \buart.Z_rx.shifter_1_LC_6_15_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_6_15_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_6_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19832),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__22069),
            .sr(N__22006));
    defparam \buart.Z_rx.shifter_fast_4_LC_6_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_6_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_6_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(bu_rx_data_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22269),
            .ce(N__22069),
            .sr(N__22006));
    defparam \uu2.w_addr_user_5_LC_7_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_7_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_7_1_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_5_LC_7_1_0  (
            .in0(N__13933),
            .in1(N__14122),
            .in2(N__14182),
            .in3(N__14207),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__14054));
    defparam \uu2.w_addr_user_4_LC_7_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_7_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_7_1_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_user_4_LC_7_1_1  (
            .in0(N__14121),
            .in1(N__13932),
            .in2(_gnd_net_),
            .in3(N__14173),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__14054));
    defparam \uu2.w_addr_user_6_LC_7_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_7_1_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_7_1_2  (
            .in0(N__13934),
            .in1(N__14123),
            .in2(N__14141),
            .in3(N__14492),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__14054));
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_7_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_7_2_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \uu2.w_addr_user_RNI93NG7_2_LC_7_2_0  (
            .in0(N__13948),
            .in1(N__15994),
            .in2(_gnd_net_),
            .in3(N__13955),
            .lcout(\uu2.un28_w_addr_user_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un20_w_addr_user_1_LC_7_2_2 .C_ON=1'b0;
    defparam \uu2.un20_w_addr_user_1_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un20_w_addr_user_1_LC_7_2_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uu2.un20_w_addr_user_1_LC_7_2_2  (
            .in0(N__13982),
            .in1(N__15854),
            .in2(N__13973),
            .in3(N__17086),
            .lcout(\uu2.un20_w_addr_userZ0Z_1 ),
            .ltout(\uu2.un20_w_addr_userZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI43E87_2_LC_7_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI43E87_2_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI43E87_2_LC_7_2_3 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \uu2.w_addr_user_RNI43E87_2_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__13949),
            .in2(N__13940),
            .in3(N__14723),
            .lcout(\uu2.w_addr_user_RNI43E87Z0Z_2 ),
            .ltout(\uu2.w_addr_user_RNI43E87Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNID65PE_2_LC_7_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNID65PE_2_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNID65PE_2_LC_7_2_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_user_RNID65PE_2_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13937),
            .in3(N__13928),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_0_LC_7_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_7_2_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_user_0_LC_7_2_5  (
            .in0(N__13929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14384),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__14047));
    defparam \uu2.w_addr_user_1_LC_7_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_7_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_user_1_LC_7_2_6  (
            .in0(N__14385),
            .in1(N__14290),
            .in2(_gnd_net_),
            .in3(N__13930),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__14047));
    defparam \uu2.w_addr_user_2_LC_7_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_7_2_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_2_LC_7_2_7  (
            .in0(N__13931),
            .in1(N__14339),
            .in2(N__14301),
            .in3(N__14386),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__14047));
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_2  (
            .in0(N__14208),
            .in1(N__14234),
            .in2(N__14464),
            .in3(N__14368),
            .lcout(\uu2.un3_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_7_3_3  (
            .in0(N__14369),
            .in1(N__14340),
            .in2(N__14244),
            .in3(N__14294),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__14069),
            .sr(N__14046));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_3_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_3_4  (
            .in0(N__14209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14181),
            .lcout(\uu2.un426_ci_3 ),
            .ltout(\uu2.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_7_3_5  (
            .in0(N__14119),
            .in1(N__14459),
            .in2(N__14144),
            .in3(N__14497),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__14069),
            .sr(N__14046));
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_7_3_6  (
            .in0(N__14134),
            .in1(N__14120),
            .in2(N__14090),
            .in3(N__14441),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__14069),
            .sr(N__14046));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_4_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_4_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_7_4_1  (
            .in0(N__15679),
            .in1(N__15986),
            .in2(N__14498),
            .in3(N__15826),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_4_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_4_2 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_7_4_2  (
            .in0(N__15827),
            .in1(N__14460),
            .in2(N__16972),
            .in3(N__15985),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_4_3 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_52_LC_7_4_3  (
            .in0(N__17256),
            .in1(N__16957),
            .in2(N__15685),
            .in3(N__16115),
            .lcout(\uu2.mem0.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI90ME1_5_LC_7_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI90ME1_5_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI90ME1_5_LC_7_4_4 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI90ME1_5_LC_7_4_4  (
            .in0(N__16114),
            .in1(N__15678),
            .in2(N__16971),
            .in3(N__17257),
            .lcout(\uu2.bitmap_pmux_sn_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_4_5 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_nesr_8_LC_7_4_5  (
            .in0(N__15680),
            .in1(N__16961),
            .in2(N__15718),
            .in3(N__16116),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_8C_net ),
            .ce(N__15611),
            .sr(N__21947));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_4_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_4_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_4_7  (
            .in0(N__14496),
            .in1(_gnd_net_),
            .in2(N__14465),
            .in3(_gnd_net_),
            .lcout(\uu2.vbuf_w_addr_user.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNILN731_40_LC_7_5_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNILN731_40_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNILN731_40_LC_7_5_0 .LUT_INIT=16'b0001100101011101;
    LogicCell40 \uu2.bitmap_RNILN731_40_LC_7_5_0  (
            .in0(N__16113),
            .in1(N__16042),
            .in2(N__14978),
            .in3(N__14435),
            .lcout(\uu2.bitmap_pmux_26_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_7_5_1 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_7_5_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_40_LC_7_5_1  (
            .in0(N__15239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20052),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__21945));
    defparam \uu2.bitmap_52_LC_7_5_2 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_7_5_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.bitmap_52_LC_7_5_2  (
            .in0(N__20053),
            .in1(_gnd_net_),
            .in2(N__14429),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__21945));
    defparam \uu2.w_addr_displaying_RNIBICU6_2_LC_7_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIBICU6_2_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIBICU6_2_LC_7_5_3 .LUT_INIT=16'b1101111111010101;
    LogicCell40 \uu2.w_addr_displaying_RNIBICU6_2_LC_7_5_3  (
            .in0(N__14411),
            .in1(N__16055),
            .in2(N__14420),
            .in3(N__14816),
            .lcout(\uu2.w_addr_displaying_RNIBICU6Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIF31A1_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIF31A1_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIF31A1_LC_7_5_4 .LUT_INIT=16'b0010101000101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNIF31A1_LC_7_5_4  (
            .in0(N__17615),
            .in1(N__17762),
            .in2(N__16126),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(\uu2.bitmap_pmux_sn_N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIBICU6_0_2_LC_7_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIBICU6_0_2_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIBICU6_0_2_LC_7_5_5 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \uu2.w_addr_displaying_RNIBICU6_0_2_LC_7_5_5  (
            .in0(N__14410),
            .in1(N__14815),
            .in2(N__14402),
            .in3(N__16054),
            .lcout(\uu2.w_addr_displaying_RNIBICU6_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIL1MV_52_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIL1MV_52_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIL1MV_52_LC_7_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.bitmap_RNIL1MV_52_LC_7_5_6  (
            .in0(N__16109),
            .in1(N__14399),
            .in2(_gnd_net_),
            .in3(N__14393),
            .lcout(),
            .ltout(\uu2.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNICS7L2_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNICS7L2_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNICS7L2_LC_7_5_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_RNICS7L2_LC_7_5_7  (
            .in0(N__17629),
            .in1(N__16949),
            .in2(N__14819),
            .in3(N__16001),
            .lcout(\uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_7_6_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_3_LC_7_6_0  (
            .in0(N__14807),
            .in1(N__14801),
            .in2(_gnd_net_),
            .in3(N__14714),
            .lcout(\Lab_UT.dictrl.un1_next_alarmstate21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sec1_1_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.sec1_1_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sec1_1_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.sec1_1_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14759),
            .lcout(\Lab_UT.sec1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI34K17_5_LC_7_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI34K17_5_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI34K17_5_LC_7_6_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_RNI34K17_5_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__14713),
            .in2(_gnd_net_),
            .in3(N__17281),
            .lcout(\uu2.N_31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_7_6_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_7_6_3 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_7_6_3  (
            .in0(N__14589),
            .in1(N__14653),
            .in2(_gnd_net_),
            .in3(N__14556),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_7_6_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_7_6_4 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_7_6_4  (
            .in0(N__14557),
            .in1(N__14591),
            .in2(N__14657),
            .in3(N__14638),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_7_6_5 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_7_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__14634),
            .in2(_gnd_net_),
            .in3(N__14651),
            .lcout(\resetGen.un241_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_7_6_6 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_7_6_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_7_6_6  (
            .in0(N__14652),
            .in1(_gnd_net_),
            .in2(N__14639),
            .in3(N__14620),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_7_6_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_7_6_7 .LUT_INIT=16'b0000000010011100;
    LogicCell40 \resetGen.reset_count_3_LC_7_6_7  (
            .in0(N__14590),
            .in1(N__14512),
            .in2(N__14561),
            .in3(N__14558),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22326),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_7_7_0 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_7_7_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_93_LC_7_7_0  (
            .in0(N__20024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18560),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \uu2.bitmap_180_LC_7_7_1 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_7_7_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_180_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__14954),
            .in2(_gnd_net_),
            .in3(N__20022),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \uu2.bitmap_111_LC_7_7_2 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_7_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14946),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \uu2.vram_rd_clk_det_0_LC_7_7_5 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_7_7_5 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_7_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14881),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \uu2.vram_rd_clk_det_1_LC_7_7_6 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_7_7_6 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_7_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14845),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \uu2.bitmap_221_LC_7_7_7 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_7_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_221_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__18599),
            .in2(_gnd_net_),
            .in3(N__20023),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__21941));
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_0_2_LC_7_8_0 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \Lab_UT.bcd2segment3.segment_0_2_LC_7_8_0  (
            .in0(N__15217),
            .in1(N__15163),
            .in2(N__15112),
            .in3(N__15024),
            .lcout(\Lab_UT.bcd2segment3.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_7_8_1 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_4_LC_7_8_1  (
            .in0(N__15158),
            .in1(N__15027),
            .in2(N__15115),
            .in3(N__15212),
            .lcout(\Lab_UT.bcd2segment3.segmentUQ_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_7_8_2 .LUT_INIT=16'b1111101111000010;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_5_LC_7_8_2  (
            .in0(N__15213),
            .in1(N__15159),
            .in2(N__15111),
            .in3(N__15023),
            .lcout(\Lab_UT.bcd2segment3.segmentUQ_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_7_8_3 .LUT_INIT=16'b1110100111100001;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_6_LC_7_8_3  (
            .in0(N__15160),
            .in1(N__15026),
            .in2(N__15114),
            .in3(N__15214),
            .lcout(\Lab_UT.bcd2segment3.segmentUQ_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_7_8_4 .LUT_INIT=16'b1101111101111001;
    LogicCell40 \Lab_UT.bcd2segment3.segment_0_0_LC_7_8_4  (
            .in0(N__15215),
            .in1(N__15161),
            .in2(N__15110),
            .in3(N__15022),
            .lcout(\Lab_UT.bcd2segment3.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segment_0_1_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_0_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_0_1_LC_7_8_5 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \Lab_UT.bcd2segment3.segment_0_1_LC_7_8_5  (
            .in0(N__15162),
            .in1(N__15028),
            .in2(N__15116),
            .in3(N__15216),
            .lcout(\Lab_UT.bcd2segment3.segment_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_7_8_6 .LUT_INIT=16'b1111100011100110;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_3_LC_7_8_6  (
            .in0(N__15218),
            .in1(N__15164),
            .in2(N__15113),
            .in3(N__15025),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_7_8_7 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_7_8_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_296_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14981),
            .in3(N__19981),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__21938));
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_9_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_7_9_0  (
            .in0(N__18464),
            .in1(N__16249),
            .in2(N__15287),
            .in3(N__15307),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_7_9_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_7_9_1  (
            .in0(N__15263),
            .in1(N__16490),
            .in2(_gnd_net_),
            .in3(N__18347),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_9_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_7_9_2  (
            .in0(N__18348),
            .in1(N__15306),
            .in2(N__14963),
            .in3(N__16248),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_7_9_3 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_7_9_3  (
            .in0(N__18525),
            .in1(N__14960),
            .in2(N__15269),
            .in3(N__19873),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_7_9_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_7_9_4  (
            .in0(N__18526),
            .in1(N__16250),
            .in2(N__15314),
            .in3(N__15308),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_9_5  (
            .in0(N__18524),
            .in1(N__18463),
            .in2(_gnd_net_),
            .in3(N__18346),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_9_6 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_9_6  (
            .in0(N__15267),
            .in1(N__19412),
            .in2(N__15311),
            .in3(N__18396),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_9_7 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_7_9_7  (
            .in0(N__15305),
            .in1(N__18397),
            .in2(N__15290),
            .in3(N__16247),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22301),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_10_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_10_0  (
            .in0(N__22760),
            .in1(N__18465),
            .in2(N__15268),
            .in3(N__18345),
            .lcout(\Lab_UT.didp.countrce1.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_4_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_4_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_4_LC_7_10_1 .LUT_INIT=16'b0100010001001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_4_LC_7_10_1  (
            .in0(N__19411),
            .in1(N__18617),
            .in2(N__19879),
            .in3(N__22759),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_0_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_0_LC_7_10_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_0_LC_7_10_2  (
            .in0(N__19138),
            .in1(N__16517),
            .in2(N__15275),
            .in3(N__19177),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_9_LC_7_10_3 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_LC_7_10_3  (
            .in0(N__19018),
            .in1(N__16508),
            .in2(N__15272),
            .in3(N__15320),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22294),
            .ce(),
            .sr(N__21979));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_8_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_8_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_8_LC_7_10_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_8_LC_7_10_4  (
            .in0(N__21753),
            .in1(N__21465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_5_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_5_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_5_LC_7_10_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_5_LC_7_10_5  (
            .in0(N__19176),
            .in1(N__23210),
            .in2(N__15242),
            .in3(N__19137),
            .lcout(\Lab_UT.dictrl.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_LC_7_10_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_LC_7_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__15392),
            .in2(_gnd_net_),
            .in3(N__19017),
            .lcout(\Lab_UT.dicLdSones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22294),
            .ce(),
            .sr(N__21979));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_6_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_6_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_6_LC_7_11_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_6_LC_7_11_0  (
            .in0(N__21063),
            .in1(N__21468),
            .in2(_gnd_net_),
            .in3(N__20828),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_4_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_4_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_4_LC_7_11_1 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_4_LC_7_11_1  (
            .in0(N__22743),
            .in1(N__19880),
            .in2(N__15338),
            .in3(N__19389),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_0_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_0_LC_7_11_2 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_0_LC_7_11_2  (
            .in0(N__16523),
            .in1(N__19140),
            .in2(N__15335),
            .in3(N__19175),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_LC_7_11_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_10_LC_7_11_3 .LUT_INIT=16'b1111111100000111;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_LC_7_11_3  (
            .in0(N__15329),
            .in1(N__16397),
            .in2(N__15332),
            .in3(N__19022),
            .lcout(\Lab_UT.LdSones_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22288),
            .ce(),
            .sr(N__21983));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_1_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_1_LC_7_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_1_LC_7_11_4  (
            .in0(N__21717),
            .in1(N__20829),
            .in2(N__20664),
            .in3(N__21469),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g3_0_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g3_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g3_0_LC_7_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g3_0_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(_gnd_net_),
            .in3(N__21062),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_7_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_7_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_7_LC_7_11_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_7_LC_7_11_6  (
            .in0(N__20395),
            .in1(N__21467),
            .in2(N__15323),
            .in3(N__23222),
            .lcout(\Lab_UT.dictrl.i6_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_1_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_1_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_1_LC_7_11_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_1_LC_7_11_7  (
            .in0(N__21470),
            .in1(N__20649),
            .in2(N__20854),
            .in3(N__21718),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_RNIOF67_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_RNIOF67_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_RNIOF67_LC_7_12_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_RNIOF67_LC_7_12_0  (
            .in0(N__21124),
            .in1(N__21427),
            .in2(N__21752),
            .in3(N__21212),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_LC_7_12_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_LC_7_12_1  (
            .in0(N__20853),
            .in1(N__15410),
            .in2(N__21763),
            .in3(N__15401),
            .lcout(\Lab_UT.dictrl.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22283),
            .ce(),
            .sr(N__21986));
    defparam \Lab_UT.dictrl.g0_1_0_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_1_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_1_0_LC_7_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.g0_1_0_LC_7_12_2  (
            .in0(N__22974),
            .in1(N__19504),
            .in2(N__20903),
            .in3(N__21572),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_8_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_8_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_8_LC_7_12_3 .LUT_INIT=16'b0001110111011101;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_8_LC_7_12_3  (
            .in0(N__20519),
            .in1(N__21125),
            .in2(N__15416),
            .in3(N__19092),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_29_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_6_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_6_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_6_LC_7_12_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_6_LC_7_12_4  (
            .in0(N__21428),
            .in1(N__21211),
            .in2(N__15413),
            .in3(N__15461),
            .lcout(\Lab_UT.dictrl.N_30_0 ),
            .ltout(\Lab_UT.dictrl.N_30_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNI6JM59_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNI6JM59_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNI6JM59_LC_7_12_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNI6JM59_LC_7_12_5  (
            .in0(N__21711),
            .in1(N__20850),
            .in2(N__15404),
            .in3(N__15400),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_2 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_RNO_0_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNO_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNO_0_LC_7_12_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNO_0_LC_7_12_6  (
            .in0(N__20851),
            .in1(N__21712),
            .in2(N__15383),
            .in3(N__18875),
            .lcout(),
            .ltout(\Lab_UT.dictrl.dicLdAMones_0_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_12_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_12_7 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_7_12_7  (
            .in0(N__21713),
            .in1(N__20852),
            .in2(N__15380),
            .in3(N__18831),
            .lcout(\Lab_UT.dicLdAMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22283),
            .ce(),
            .sr(N__21986));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_13_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_13_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_13_LC_7_13_0 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_13_LC_7_13_0  (
            .in0(N__22531),
            .in1(N__19460),
            .in2(N__15362),
            .in3(N__19256),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_LC_7_13_1 .LUT_INIT=16'b0101001111001110;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_LC_7_13_1  (
            .in0(N__23209),
            .in1(N__21109),
            .in2(N__15500),
            .in3(N__16727),
            .lcout(\Lab_UT.dictrl.N_7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_5_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_5_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_5_LC_7_13_2 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_5_LC_7_13_2  (
            .in0(N__16664),
            .in1(N__19592),
            .in2(N__15527),
            .in3(N__19541),
            .lcout(\Lab_UT.dictrl.g2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_1_2_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_1_2_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_1_2_LC_7_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_1_2_LC_7_13_3  (
            .in0(N__19540),
            .in1(N__16663),
            .in2(N__15491),
            .in3(N__16711),
            .lcout(\Lab_UT.dictrl.g0_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_4_2_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_4_2_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_4_2_LC_7_13_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.g0_4_2_LC_7_13_4  (
            .in0(N__16712),
            .in1(N__19593),
            .in2(N__16670),
            .in3(N__19542),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_10_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_10_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_10_LC_7_13_5 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \Lab_UT.dictrl.g0_10_LC_7_13_5  (
            .in0(N__21569),
            .in1(N__20494),
            .in2(N__15473),
            .in3(N__22969),
            .lcout(\Lab_UT.dictrl.next_state18_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_LC_7_13_6 .LUT_INIT=16'b0101010101011111;
    LogicCell40 \Lab_UT.dictrl.g1_0_LC_7_13_6  (
            .in0(N__22970),
            .in1(_gnd_net_),
            .in2(N__20498),
            .in3(N__21570),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_LC_7_13_7 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_1_LC_7_13_7  (
            .in0(N__18890),
            .in1(N__22532),
            .in2(N__15464),
            .in3(N__21110),
            .lcout(\Lab_UT.dictrl.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_2_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_2_LC_7_14_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_2_LC_7_14_0  (
            .in0(N__19545),
            .in1(N__16659),
            .in2(N__19600),
            .in3(N__16715),
            .lcout(\Lab_UT.dictrl.next_state12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_2_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_2_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_2_LC_7_14_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_1_2_LC_7_14_1  (
            .in0(N__16714),
            .in1(N__19588),
            .in2(N__16668),
            .in3(N__19544),
            .lcout(\Lab_UT.dictrl.g2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state32_4_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state32_4_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state32_4_LC_7_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.next_state32_4_LC_7_14_2  (
            .in0(N__19543),
            .in1(N__16655),
            .in2(N__19599),
            .in3(N__16713),
            .lcout(\Lab_UT.dictrl.next_state32Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_5_LC_7_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_7_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_7_14_4  (
            .in0(N__22870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22274),
            .ce(N__22068),
            .sr(N__22007));
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_rep1_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_rep1_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22869),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22274),
            .ce(N__22068),
            .sr(N__22007));
    defparam \buart.Z_rx.shifter_4_rep1_LC_7_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep1_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_rep1_LC_7_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_rep1_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22545),
            .lcout(bu_rx_data_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22274),
            .ce(N__22068),
            .sr(N__22007));
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23034),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22271),
            .ce(N__22067),
            .sr(N__22008));
    defparam \buart.Z_rx.shifter_fast_3_LC_7_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_7_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22458),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22271),
            .ce(N__22067),
            .sr(N__22008));
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_3_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_45_LC_8_3_0  (
            .in0(N__17507),
            .in1(N__17888),
            .in2(_gnd_net_),
            .in3(N__17631),
            .lcout(\uu2.mem0.G_11_0_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_3_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_8_3_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_53_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__17506),
            .in2(_gnd_net_),
            .in3(N__17758),
            .lcout(),
            .ltout(\uu2.mem0.N_98_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_3_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_8_3_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_46_LC_8_3_2  (
            .in0(N__17990),
            .in1(N__17632),
            .in2(N__15512),
            .in3(N__17551),
            .lcout(),
            .ltout(\uu2.mem0.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_3_3 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_30_LC_8_3_3  (
            .in0(N__15509),
            .in1(N__17202),
            .in2(N__15503),
            .in3(N__17420),
            .lcout(),
            .ltout(\uu2.mem0.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_8_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_8_3_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_20_LC_8_3_4  (
            .in0(N__15587),
            .in1(N__17119),
            .in2(N__15578),
            .in3(N__16785),
            .lcout(\uu2.mem0.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_8_3_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_8_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_23_LC_8_3_5  (
            .in0(N__15671),
            .in1(N__16962),
            .in2(N__18117),
            .in3(N__16119),
            .lcout(\uu2.mem0.G_11_0_0_a2_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_8_3_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_28_LC_8_3_6  (
            .in0(N__16120),
            .in1(_gnd_net_),
            .in2(N__16973),
            .in3(_gnd_net_),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI31F32_34_LC_8_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI31F32_34_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI31F32_34_LC_8_4_0 .LUT_INIT=16'b0000110011111010;
    LogicCell40 \uu2.bitmap_RNI31F32_34_LC_8_4_0  (
            .in0(N__19922),
            .in1(N__19673),
            .in2(N__17633),
            .in3(N__15575),
            .lcout(),
            .ltout(\uu2.bitmap_RNI31F32Z0Z_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNII6975_34_LC_8_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNII6975_34_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNII6975_34_LC_8_4_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.bitmap_RNII6975_34_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__15533),
            .in2(N__15569),
            .in3(N__15539),
            .lcout(),
            .ltout(\uu2.N_401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI8B24J_34_LC_8_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI8B24J_34_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI8B24J_34_LC_8_4_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \uu2.bitmap_RNI8B24J_34_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__15566),
            .in2(N__15560),
            .in3(N__15557),
            .lcout(\uu2.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIJS4P_162_LC_8_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJS4P_162_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJS4P_162_LC_8_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIJS4P_162_LC_8_4_3  (
            .in0(N__16041),
            .in1(N__16190),
            .in2(_gnd_net_),
            .in3(N__19664),
            .lcout(),
            .ltout(\uu2.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_8_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_8_4_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uu2.bitmap_RNI2Q8F1_111_LC_8_4_4  (
            .in0(N__15551),
            .in1(_gnd_net_),
            .in2(N__15542),
            .in3(N__15623),
            .lcout(\uu2.bitmap_RNI2Q8F1Z0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIDBHK1_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIDBHK1_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIDBHK1_LC_8_4_5 .LUT_INIT=16'b0000000001110110;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNIDBHK1_LC_8_4_5  (
            .in0(N__17741),
            .in1(N__17541),
            .in2(N__17630),
            .in3(N__16950),
            .lcout(\uu2.bitmap_pmux_sn_N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_8_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_8_4_6 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_8_4_6  (
            .in0(N__15617),
            .in1(N__16040),
            .in2(_gnd_net_),
            .in3(N__17332),
            .lcout(\uu2.bitmap_pmux_sn_N_54_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_8_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_8_5_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_3_LC_8_5_0  (
            .in0(N__17389),
            .in1(N__17205),
            .in2(N__16046),
            .in3(N__17884),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_8_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_8_5_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_LC_8_5_1  (
            .in0(N__17203),
            .in1(N__17628),
            .in2(N__17910),
            .in3(N__17390),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.w_addr_displaying_nesr_1_LC_8_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_1_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_1_LC_8_5_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_nesr_1_LC_8_5_2  (
            .in0(N__17988),
            .in1(_gnd_net_),
            .in2(N__17764),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_8_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_8_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__17750),
            .in2(_gnd_net_),
            .in3(N__17986),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.w_addr_displaying_nesr_3_LC_8_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_8_5_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_8_5_5  (
            .in0(N__17204),
            .in1(N__18072),
            .in2(N__17911),
            .in3(N__17391),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_8_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_8_5_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_1_LC_8_5_6  (
            .in0(N__17987),
            .in1(_gnd_net_),
            .in2(N__17763),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_3C_net ),
            .ce(N__15607),
            .sr(N__21948));
    defparam \uu2.bitmap_RNIFH0N_90_LC_8_6_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIFH0N_90_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIFH0N_90_LC_8_6_0 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \uu2.bitmap_RNIFH0N_90_LC_8_6_0  (
            .in0(N__18308),
            .in1(N__18179),
            .in2(N__18236),
            .in3(N__15593),
            .lcout(\uu2.bitmap_pmux_19_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_90_LC_8_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_8_6_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_90_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__18587),
            .in2(_gnd_net_),
            .in3(N__20021),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__21946));
    defparam \uu2.bitmap_186_LC_8_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_8_6_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_186_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__18578),
            .in2(_gnd_net_),
            .in3(N__20019),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__21946));
    defparam \uu2.bitmap_RNIKGSI_58_LC_8_6_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKGSI_58_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKGSI_58_LC_8_6_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNIKGSI_58_LC_8_6_4  (
            .in0(N__16169),
            .in1(N__18180),
            .in2(_gnd_net_),
            .in3(N__16133),
            .lcout(),
            .ltout(\uu2.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI04AD1_314_LC_8_6_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI04AD1_314_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI04AD1_314_LC_8_6_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.bitmap_RNI04AD1_314_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__16125),
            .in2(N__16058),
            .in3(N__16010),
            .lcout(\uu2.bitmap_RNI04AD1Z0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_314_LC_8_6_6 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_8_6_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_314_LC_8_6_6  (
            .in0(N__20020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18608),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__21946));
    defparam \uu2.bitmap_RNICM7R_180_LC_8_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNICM7R_180_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNICM7R_180_LC_8_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.bitmap_RNICM7R_180_LC_8_6_7  (
            .in0(N__16039),
            .in1(N__16016),
            .in2(_gnd_net_),
            .in3(N__16009),
            .lcout(\uu2.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_7_LC_8_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_7_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_8_7_3  (
            .in0(N__17297),
            .in1(N__15657),
            .in2(N__18188),
            .in3(N__15724),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_7C_net ),
            .ce(),
            .sr(N__21944));
    defparam \uu2.w_addr_displaying_7_LC_8_7_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_8_7_5 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \uu2.w_addr_displaying_7_LC_8_7_5  (
            .in0(N__17296),
            .in1(N__15656),
            .in2(N__16966),
            .in3(N__15723),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_7C_net ),
            .ce(),
            .sr(N__21944));
    defparam \uu2.w_addr_displaying_RNIVAPV6_5_LC_8_7_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIVAPV6_5_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIVAPV6_5_LC_8_7_6 .LUT_INIT=16'b1111111101011101;
    LogicCell40 \uu2.w_addr_displaying_RNIVAPV6_5_LC_8_7_6  (
            .in0(N__15929),
            .in1(N__15754),
            .in2(N__15725),
            .in3(N__15855),
            .lcout(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5 ),
            .ltout(\uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_6_LC_8_7_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_LC_8_7_7 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_LC_8_7_7 .LUT_INIT=16'b1110111110110000;
    LogicCell40 \uu2.w_addr_displaying_6_LC_8_7_7  (
            .in0(N__15755),
            .in1(N__15722),
            .in2(N__15692),
            .in3(N__15658),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_7C_net ),
            .ce(),
            .sr(N__21944));
    defparam \uu2.bitmap_203_LC_8_8_0 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_8_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_203_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__16208),
            .in2(_gnd_net_),
            .in3(N__19976),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \uu2.bitmap_200_LC_8_8_1 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_8_8_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_200_LC_8_8_1  (
            .in0(N__19975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16202),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \uu2.bitmap_168_LC_8_8_2 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_8_8_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_168_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__16196),
            .in2(_gnd_net_),
            .in3(N__19974),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \uu2.bitmap_75_LC_8_8_3 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_8_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_75_LC_8_8_3  (
            .in0(N__19979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16181),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \uu2.bitmap_72_LC_8_8_4 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_8_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_72_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__16175),
            .in2(_gnd_net_),
            .in3(N__19978),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \uu2.bitmap_58_LC_8_8_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_8_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_58_LC_8_8_5  (
            .in0(N__19977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18566),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__21939));
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_9_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_9_0 .LUT_INIT=16'b1011101110101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_LC_8_9_0  (
            .in0(N__20848),
            .in1(N__21269),
            .in2(N__19043),
            .in3(N__21740),
            .lcout(\Lab_UT.state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22310),
            .ce(),
            .sr(N__21980));
    defparam \Lab_UT.dictrl.state_ret_5_RNIIMGL_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_RNIIMGL_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_RNIIMGL_LC_8_9_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_RNIIMGL_LC_8_9_1  (
            .in0(N__21738),
            .in1(N__18805),
            .in2(_gnd_net_),
            .in3(N__23181),
            .lcout(\Lab_UT.LdASones ),
            .ltout(\Lab_UT.LdASones_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNO_0_0_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNO_0_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNO_0_0_LC_8_9_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Lab_UT.didp.ce_RNO_0_0_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16148),
            .in3(N__16145),
            .lcout(\Lab_UT.didp.ce_9_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_RNI0TGF_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_RNI0TGF_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_RNI0TGF_LC_8_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_RNI0TGF_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__18670),
            .in2(_gnd_net_),
            .in3(N__20606),
            .lcout(\Lab_UT.dicRun_2 ),
            .ltout(\Lab_UT.dicRun_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_0_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_8_9_4 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \Lab_UT.didp.ce_0_LC_8_9_4  (
            .in0(N__18806),
            .in1(N__16355),
            .in2(N__16349),
            .in3(N__16334),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22310),
            .ce(),
            .sr(N__21980));
    defparam \Lab_UT.dictrl.state_ret_1_RNIKRKU_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_RNIKRKU_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_RNIKRKU_LC_8_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_RNIKRKU_LC_8_9_5  (
            .in0(N__18804),
            .in1(N__20605),
            .in2(_gnd_net_),
            .in3(N__18669),
            .lcout(\Lab_UT.Run ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_9_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_9_6 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_LC_8_9_6  (
            .in0(N__20849),
            .in1(N__21739),
            .in2(N__20534),
            .in3(N__16538),
            .lcout(\Lab_UT.dictrl.state_i_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22310),
            .ce(),
            .sr(N__21980));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_3_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_3_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_3_LC_8_10_0 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_3_LC_8_10_0  (
            .in0(N__19352),
            .in1(N__22765),
            .in2(N__19871),
            .in3(N__16220),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_0_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_0_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_0_LC_8_10_1 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_0_LC_8_10_1  (
            .in0(N__16214),
            .in1(N__16229),
            .in2(N__16223),
            .in3(N__18772),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_LC_8_10_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_LC_8_10_2  (
            .in0(N__20811),
            .in1(N__18878),
            .in2(N__21794),
            .in3(N__18838),
            .lcout(\Lab_UT.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22302),
            .ce(),
            .sr(N__21984));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_7_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_7_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_7_LC_8_10_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_7_LC_8_10_3  (
            .in0(N__20795),
            .in1(N__21064),
            .in2(_gnd_net_),
            .in3(N__16593),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_4_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_4_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_4_LC_8_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_4_LC_8_10_4  (
            .in0(N__21784),
            .in1(N__21369),
            .in2(_gnd_net_),
            .in3(N__23203),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_3_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_3_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_3_LC_8_10_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_3_LC_8_10_5  (
            .in0(N__23204),
            .in1(N__21786),
            .in2(_gnd_net_),
            .in3(N__16594),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_3_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_3_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_3_LC_8_10_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_3_LC_8_10_7  (
            .in0(N__23205),
            .in1(N__21785),
            .in2(_gnd_net_),
            .in3(N__16595),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_2_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_2_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_2_LC_8_11_0 .LUT_INIT=16'b1011101110110001;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_2_LC_8_11_0  (
            .in0(N__21060),
            .in1(N__19201),
            .in2(N__16622),
            .in3(N__18773),
            .lcout(\Lab_UT.dictrl.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_7_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_7_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_7_LC_8_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_7_LC_8_11_1  (
            .in0(N__20817),
            .in1(N__21059),
            .in2(_gnd_net_),
            .in3(N__16591),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_3_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_3_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_3_LC_8_11_2 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_3_LC_8_11_2  (
            .in0(N__19338),
            .in1(N__19833),
            .in2(N__16496),
            .in3(N__22741),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_8_11_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_LC_8_11_3  (
            .in0(N__16760),
            .in1(N__16751),
            .in2(N__22875),
            .in3(N__16482),
            .lcout(\Lab_UT.dictrl.next_alarmstateZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m4_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m4_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m4_LC_8_11_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m4_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__23192),
            .in2(_gnd_net_),
            .in3(N__20394),
            .lcout(\Lab_UT.dictrl.N_5 ),
            .ltout(\Lab_UT.dictrl.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_2_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_2_LC_8_11_5 .LUT_INIT=16'b1111101000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_2_LC_8_11_5  (
            .in0(N__16604),
            .in1(N__19200),
            .in2(N__16400),
            .in3(N__21061),
            .lcout(\Lab_UT.dictrl.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_5_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_5_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_5_LC_8_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_5_LC_8_11_6  (
            .in0(N__16610),
            .in1(N__19139),
            .in2(N__19178),
            .in3(N__23193),
            .lcout(\Lab_UT.dictrl.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_5_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_5_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_5_LC_8_11_7 .LUT_INIT=16'b1100100011111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_5_LC_8_11_7  (
            .in0(N__22742),
            .in1(N__19339),
            .in2(N__19870),
            .in3(N__16592),
            .lcout(\Lab_UT.dictrl.g0_0_0_o4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_1_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_1_LC_8_12_0 .LUT_INIT=16'b0001111100000000;
    LogicCell40 \Lab_UT.dictrl.g0_1_LC_8_12_0  (
            .in0(N__19503),
            .in1(N__16860),
            .in2(N__22975),
            .in3(N__16576),
            .lcout(\Lab_UT.dictrl.next_state18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_11_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_11_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_11_LC_8_12_1 .LUT_INIT=16'b0101010011111110;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_11_LC_8_12_1  (
            .in0(N__21209),
            .in1(N__19184),
            .in2(N__21485),
            .in3(N__16681),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_10_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_10_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_10_LC_8_12_2 .LUT_INIT=16'b1010111100100111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_10_LC_8_12_2  (
            .in0(N__21111),
            .in1(N__16556),
            .in2(N__16613),
            .in3(N__18770),
            .lcout(\Lab_UT.dictrl.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_8_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_8_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_8_LC_8_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_8_LC_8_12_3  (
            .in0(N__21431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21693),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_RNO_5_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_5_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_RNO_5_LC_8_12_4 .LUT_INIT=16'b1100100011111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_RNO_5_LC_8_12_4  (
            .in0(N__22747),
            .in1(N__19364),
            .in2(N__19855),
            .in3(N__16578),
            .lcout(\Lab_UT.dictrl.g0_0_i_o4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_4_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_4_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_4_LC_8_12_5 .LUT_INIT=16'b0000001010101010;
    LogicCell40 \Lab_UT.dictrl.g0_4_LC_8_12_5  (
            .in0(N__16577),
            .in1(N__21555),
            .in2(N__20493),
            .in3(N__22965),
            .lcout(\Lab_UT.dictrl.next_state18_0 ),
            .ltout(\Lab_UT.dictrl.next_state18_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_3_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_3_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_3_LC_8_12_6 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_3_LC_8_12_6  (
            .in0(N__16682),
            .in1(_gnd_net_),
            .in2(N__16550),
            .in3(N__21112),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_9_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_9_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_9_LC_8_12_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_9_LC_8_12_7  (
            .in0(N__21432),
            .in1(N__20645),
            .in2(N__16547),
            .in3(N__16544),
            .lcout(\Lab_UT.dictrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_13_0 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_13_0  (
            .in0(N__21530),
            .in1(N__20460),
            .in2(N__22971),
            .in3(N__16529),
            .lcout(\Lab_UT.dictrl.g2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_LC_8_13_1 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g1_LC_8_13_1  (
            .in0(N__19707),
            .in1(N__19453),
            .in2(_gnd_net_),
            .in3(N__19249),
            .lcout(\Lab_UT.dictrl.gZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_3_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_3_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_3_LC_8_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_3_LC_8_13_2  (
            .in0(N__16862),
            .in1(N__22455),
            .in2(N__19505),
            .in3(N__19556),
            .lcout(\Lab_UT.dictrl.next_alarmstate4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_8_13_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_0_LC_8_13_3  (
            .in0(N__19708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16716),
            .lcout(\Lab_UT.dictrl.next_alarmstate4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_0_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_0_LC_8_13_4 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_0_LC_8_13_4  (
            .in0(N__16742),
            .in1(N__22952),
            .in2(N__21554),
            .in3(N__20461),
            .lcout(\Lab_UT.dictrl.g2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_3_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_3_LC_8_13_5 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_3_LC_8_13_5  (
            .in0(N__16669),
            .in1(N__16861),
            .in2(N__19712),
            .in3(N__16717),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_0_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_0_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_0_LC_8_13_6 .LUT_INIT=16'b0000000110101011;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_1_0_LC_8_13_6  (
            .in0(N__21108),
            .in1(N__19511),
            .in2(N__16736),
            .in3(N__16733),
            .lcout(\Lab_UT.dictrl.g0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_6_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_6_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_6_LC_8_14_0 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \Lab_UT.dictrl.g0_6_LC_8_14_0  (
            .in0(N__19452),
            .in1(N__19594),
            .in2(N__19699),
            .in3(N__19248),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_LC_8_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_LC_8_14_1  (
            .in0(N__23046),
            .in1(N__22865),
            .in2(N__16721),
            .in3(N__16718),
            .lcout(\Lab_UT.dictrl.next_state12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_8_3_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_8_3_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_8_3_LC_8_14_2 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.dictrl.g0_8_3_LC_8_14_2  (
            .in0(N__19451),
            .in1(N__16654),
            .in2(N__19698),
            .in3(N__19247),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_8Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_8_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_8_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_8_LC_8_14_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_8_LC_8_14_3  (
            .in0(N__23045),
            .in1(N__22430),
            .in2(N__16877),
            .in3(N__22544),
            .lcout(\Lab_UT.dictrl.next_state12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_3_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_3_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_1_3_LC_8_14_4 .LUT_INIT=16'b1110101011111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_1_3_LC_8_14_4  (
            .in0(N__19694),
            .in1(N__16859),
            .in2(N__19499),
            .in3(N__19595),
            .lcout(\Lab_UT.dictrl.g2_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep1_LC_8_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19780),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22275),
            .ce(N__22070),
            .sr(N__22009));
    defparam \buart.Z_rx.shifter_3_LC_8_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_8_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22457),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22275),
            .ce(N__22070),
            .sr(N__22009));
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_9_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_9_3_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_18_LC_9_3_0  (
            .in0(N__16838),
            .in1(N__16810),
            .in2(N__17120),
            .in3(N__17570),
            .lcout(),
            .ltout(\uu2.mem0.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_9_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_9_3_1  (
            .in0(N__16832),
            .in1(N__17057),
            .in2(N__16826),
            .in3(N__16766),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_9_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_9_3_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__17757),
            .in2(_gnd_net_),
            .in3(N__17989),
            .lcout(\uu2.N_30_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_9_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_9_3_4 .LUT_INIT=16'b0010110110110100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_32_LC_9_3_4  (
            .in0(N__17514),
            .in1(N__18102),
            .in2(N__17207),
            .in3(N__17419),
            .lcout(),
            .ltout(\uu2.mem0.N_24_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_9_3_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_9_3_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_22_LC_9_3_5  (
            .in0(N__16811),
            .in1(N__17118),
            .in2(N__16790),
            .in3(N__16786),
            .lcout(\uu2.mem0.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_9_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_9_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_24_LC_9_3_6  (
            .in0(N__17513),
            .in1(N__17261),
            .in2(N__17206),
            .in3(N__18288),
            .lcout(),
            .ltout(\uu2.mem0.G_11_0_0_a2_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_9_3_7 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_9_3_7  (
            .in0(N__17126),
            .in1(N__17117),
            .in2(N__17093),
            .in3(N__17090),
            .lcout(\uu2.mem0.G_11_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_9_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_9_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_87_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__17051),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__21952));
    defparam \uu2.bitmap_84_LC_9_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_9_4_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_84_LC_9_4_1  (
            .in0(N__20056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17039),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__21952));
    defparam \uu2.bitmap_212_LC_9_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_9_4_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_212_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__17027),
            .in2(_gnd_net_),
            .in3(N__20054),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__21952));
    defparam \uu2.bitmap_215_LC_9_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_9_4_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_215_LC_9_4_3  (
            .in0(N__20055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17015),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__21952));
    defparam \uu2.bitmap_RNIOPSS_212_LC_9_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIOPSS_212_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIOPSS_212_LC_9_4_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \uu2.bitmap_RNIOPSS_212_LC_9_4_4  (
            .in0(N__17003),
            .in1(N__18187),
            .in2(N__16997),
            .in3(N__18226),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_17_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIEMII1_84_LC_9_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIEMII1_84_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIEMII1_84_LC_9_4_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \uu2.bitmap_RNIEMII1_84_LC_9_4_5  (
            .in0(N__16988),
            .in1(N__16982),
            .in2(N__16976),
            .in3(N__16967),
            .lcout(\uu2.N_104 ),
            .ltout(\uu2.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_9_4_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_9_4_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_38_LC_9_4_6  (
            .in0(N__18284),
            .in1(N__17627),
            .in2(N__17576),
            .in3(N__17681),
            .lcout(),
            .ltout(\uu2.mem0.G_11_0_0_a3_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_4_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_9_4_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_27_LC_9_4_7  (
            .in0(N__17435),
            .in1(N__17564),
            .in2(N__17573),
            .in3(N__18260),
            .lcout(\uu2.mem0.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_9_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_9_5_0 .LUT_INIT=16'b0100001000100001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_40_LC_9_5_0  (
            .in0(N__17387),
            .in1(N__17545),
            .in2(N__17889),
            .in3(N__17515),
            .lcout(\uu2.mem0.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_5_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_LC_9_5_1  (
            .in0(N__17547),
            .in1(N__17303),
            .in2(N__17418),
            .in3(N__17865),
            .lcout(\uu2.w_addr_displaying_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__21950));
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_9_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_9_5_2 .LUT_INIT=16'b1000010001000010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_41_LC_9_5_2  (
            .in0(N__17749),
            .in1(N__17546),
            .in2(N__17890),
            .in3(N__17516),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_9_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_9_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__17864),
            .in2(_gnd_net_),
            .in3(N__17298),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__21950));
    defparam \uu2.w_addr_displaying_fast_2_LC_9_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_9_5_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_9_5_4  (
            .in0(N__17388),
            .in1(N__17880),
            .in2(N__17315),
            .in3(N__17333),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__21950));
    defparam \uu2.w_addr_displaying_fast_0_LC_9_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__17302),
            .in2(_gnd_net_),
            .in3(N__18235),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__21950));
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_5_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_9_5_6  (
            .in0(N__17977),
            .in1(_gnd_net_),
            .in2(N__17314),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__21950));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_0_LC_9_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_0_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_0_LC_9_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_0_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__17748),
            .in2(_gnd_net_),
            .in3(N__17976),
            .lcout(\uu2.N_30_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_194_LC_9_6_0 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_9_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_194_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__19646),
            .in2(_gnd_net_),
            .in3(N__20030),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__21949));
    defparam \uu2.bitmap_66_LC_9_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_9_6_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_66_LC_9_6_1  (
            .in0(N__20032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19637),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__21949));
    defparam \uu2.bitmap_RNILQ2M_66_LC_9_6_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNILQ2M_66_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNILQ2M_66_LC_9_6_2 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \uu2.bitmap_RNILQ2M_66_LC_9_6_2  (
            .in0(N__18241),
            .in1(N__18183),
            .in2(N__17699),
            .in3(N__17690),
            .lcout(\uu2.bitmap_pmux_20_ns_1 ),
            .ltout(\uu2.bitmap_pmux_20_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_9_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_9_6_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_48_LC_9_6_3  (
            .in0(N__17662),
            .in1(N__17671),
            .in2(N__17684),
            .in3(N__17985),
            .lcout(\uu2.mem0.N_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_197_LC_9_6_4 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_9_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_197_LC_9_6_4  (
            .in0(N__19655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20031),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__21949));
    defparam \uu2.bitmap_69_LC_9_6_5 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_9_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_69_LC_9_6_5  (
            .in0(N__20033),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20354),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__21949));
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_9_6_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_9_6_6 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_33_LC_9_6_6  (
            .in0(N__17672),
            .in1(N__17663),
            .in2(N__17904),
            .in3(N__17654),
            .lcout(),
            .ltout(\uu2.mem0.N_108_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_9_6_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_9_6_7 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_25_LC_9_6_7  (
            .in0(N__18025),
            .in1(N__17771),
            .in2(N__17648),
            .in3(N__17999),
            .lcout(\uu2.mem0.N_404_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_9_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_9_7_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_55_LC_9_7_0  (
            .in0(N__18182),
            .in1(N__18251),
            .in2(N__18242),
            .in3(N__18196),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_16_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_9_7_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_49_LC_9_7_1  (
            .in0(N__18145),
            .in1(N__18130),
            .in2(N__18299),
            .in3(N__17991),
            .lcout(),
            .ltout(\uu2.mem0.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_9_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_9_7_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_39_LC_9_7_2  (
            .in0(N__18292),
            .in1(N__18114),
            .in2(N__18263),
            .in3(N__17936),
            .lcout(\uu2.mem0.G_11_0_0_a3_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_7_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_7_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_54_LC_9_7_3  (
            .in0(N__18250),
            .in1(N__18237),
            .in2(N__18200),
            .in3(N__18181),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_9_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_9_7_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_47_LC_9_7_4  (
            .in0(N__17992),
            .in1(N__18146),
            .in2(N__18134),
            .in3(N__18131),
            .lcout(),
            .ltout(\uu2.mem0.N_22_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_9_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_9_7_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_35_LC_9_7_5  (
            .in0(N__18115),
            .in1(N__18026),
            .in2(N__18011),
            .in3(N__18008),
            .lcout(\uu2.mem0.bitmap_pmux_27_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_9_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_9_7_6 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_50_LC_9_7_6  (
            .in0(N__17993),
            .in1(N__17800),
            .in2(N__17786),
            .in3(N__17929),
            .lcout(\uu2.mem0.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_9_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_9_7_7 .LUT_INIT=16'b1101010110010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_34_LC_9_7_7  (
            .in0(N__17930),
            .in1(N__17903),
            .in2(N__17804),
            .in3(N__17785),
            .lcout(\uu2.mem0.N_109_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_8_0 .LUT_INIT=16'b1111100111100010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_8_0  (
            .in0(N__18546),
            .in1(N__18482),
            .in2(N__18429),
            .in3(N__18369),
            .lcout(\Lab_UT.bcd2segment1.segmentUQ_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_9_8_1 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_2_LC_9_8_1  (
            .in0(N__18366),
            .in1(N__18414),
            .in2(N__18497),
            .in3(N__18543),
            .lcout(\Lab_UT.bcd2segment1.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_9_8_2 .LUT_INIT=16'b1110110111100100;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_5_LC_9_8_2  (
            .in0(N__18545),
            .in1(N__18483),
            .in2(N__18428),
            .in3(N__18368),
            .lcout(\Lab_UT.bcd2segment1.segmentUQ_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_9_8_3 .LUT_INIT=16'b1110110011000011;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_6_LC_9_8_3  (
            .in0(N__18365),
            .in1(N__18413),
            .in2(N__18495),
            .in3(N__18542),
            .lcout(\Lab_UT.bcd2segment1.segmentUQ_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_9_8_4 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_0_LC_9_8_4  (
            .in0(N__18547),
            .in1(N__18487),
            .in2(N__18430),
            .in3(N__18370),
            .lcout(\Lab_UT.bcd2segment1.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_0_1_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_1_LC_9_8_5 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_1_LC_9_8_5  (
            .in0(N__18367),
            .in1(N__18415),
            .in2(N__18496),
            .in3(N__18544),
            .lcout(\Lab_UT.bcd2segment1.segment_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_9_8_6 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_4_LC_9_8_6  (
            .in0(N__18548),
            .in1(N__18494),
            .in2(N__18431),
            .in3(N__18371),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_218_LC_9_8_7 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_9_8_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_218_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18311),
            .in3(N__19980),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_218C_net ),
            .ce(),
            .sr(N__21942));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_6_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_6_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_6_LC_9_9_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_6_LC_9_9_0  (
            .in0(N__18968),
            .in1(N__21374),
            .in2(_gnd_net_),
            .in3(N__20951),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_2_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_2_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_2_LC_9_9_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_2_LC_9_9_1  (
            .in0(N__21376),
            .in1(N__19208),
            .in2(N__18734),
            .in3(N__21073),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_LC_9_9_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_7_LC_9_9_2 .LUT_INIT=16'b1111111100010011;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_LC_9_9_2  (
            .in0(N__20741),
            .in1(N__18731),
            .in2(N__18725),
            .in3(N__19013),
            .lcout(\Lab_UT.LdStens_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__21985));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m33_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m33_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m33_LC_9_9_3 .LUT_INIT=16'b0100110000001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m33_LC_9_9_3  (
            .in0(N__20952),
            .in1(N__20608),
            .in2(N__21423),
            .in3(N__18969),
            .lcout(\Lab_UT.dictrl.N_39_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_6_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_6_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_6_LC_9_9_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_6_LC_9_9_4  (
            .in0(N__18967),
            .in1(N__21373),
            .in2(_gnd_net_),
            .in3(N__20950),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_2_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_2_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_2_LC_9_9_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_2_LC_9_9_5  (
            .in0(N__21375),
            .in1(N__19207),
            .in2(N__18722),
            .in3(N__21072),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_LC_9_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_6_LC_9_9_6 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_LC_9_9_6  (
            .in0(N__20876),
            .in1(N__18743),
            .in2(N__18719),
            .in3(N__19012),
            .lcout(\Lab_UT.LdStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(),
            .sr(N__21985));
    defparam \Lab_UT.didp.ce_10_1_LC_9_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_10_1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_10_1_LC_9_9_7 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \Lab_UT.didp.ce_10_1_LC_9_9_7  (
            .in0(N__20728),
            .in1(N__18671),
            .in2(N__18656),
            .in3(N__20607),
            .lcout(\Lab_UT.didp.ce_10_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m27_LC_9_10_0 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m27_LC_9_10_0  (
            .in0(N__21067),
            .in1(N__21448),
            .in2(N__21236),
            .in3(N__18632),
            .lcout(\Lab_UT.dictrl.i6_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNO_6_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_6_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNO_6_LC_9_10_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNO_6_LC_9_10_1  (
            .in0(N__21446),
            .in1(N__20796),
            .in2(_gnd_net_),
            .in3(N__21065),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m18_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m18_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m18_LC_9_10_2 .LUT_INIT=16'b1000110110101111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m18_LC_9_10_2  (
            .in0(N__21066),
            .in1(N__18769),
            .in2(N__21235),
            .in3(N__21601),
            .lcout(\Lab_UT.dictrl.N_19 ),
            .ltout(\Lab_UT.dictrl.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNICIPPD_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNICIPPD_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNICIPPD_LC_9_10_3 .LUT_INIT=16'b0000000100100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNICIPPD_LC_9_10_3  (
            .in0(N__21447),
            .in1(N__20797),
            .in2(N__18851),
            .in3(N__21619),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_RNO_1_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_RNO_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_RNO_1_LC_9_10_4 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_RNO_1_LC_9_10_4  (
            .in0(N__20798),
            .in1(N__21793),
            .in2(N__18848),
            .in3(N__18876),
            .lcout(\Lab_UT.dictrl.state_ret_5_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_LC_9_10_5 .LUT_INIT=16'b0000000100110000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_LC_9_10_5  (
            .in0(N__18845),
            .in1(N__20800),
            .in2(N__21466),
            .in3(N__21620),
            .lcout(\Lab_UT.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22311),
            .ce(),
            .sr(N__21987));
    defparam \Lab_UT.dictrl.state_ret_5_RNO_0_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_RNO_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_RNO_0_LC_9_10_6 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_RNO_0_LC_9_10_6  (
            .in0(N__20799),
            .in1(N__18877),
            .in2(N__21792),
            .in3(N__19005),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_LC_9_10_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_LC_9_10_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__18839),
            .in2(N__18815),
            .in3(N__18812),
            .lcout(\Lab_UT.dicRun_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22311),
            .ce(),
            .sr(N__21987));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_4_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_4_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_4_LC_9_11_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_4_LC_9_11_0  (
            .in0(N__21777),
            .in1(N__21364),
            .in2(_gnd_net_),
            .in3(N__23195),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_0_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_0_LC_9_11_1 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_0_LC_9_11_1  (
            .in0(N__18791),
            .in1(N__18782),
            .in2(N__18776),
            .in3(N__18771),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_9_11_2 .LUT_INIT=16'b0100010011000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_2_LC_9_11_2  (
            .in0(N__21377),
            .in1(N__19036),
            .in2(N__18977),
            .in3(N__20943),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_15_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_12_LC_9_11_3 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_LC_9_11_3  (
            .in0(N__19892),
            .in1(N__18896),
            .in2(N__19025),
            .in3(N__19011),
            .lcout(\Lab_UT.dictrl.un1_next_state66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22303),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_RNITITL_LC_9_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_RNITITL_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_RNITITL_LC_9_11_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_RNITITL_LC_9_11_4  (
            .in0(N__21776),
            .in1(N__21363),
            .in2(N__18976),
            .in3(N__23194),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_9_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_9_11_5 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_4_LC_9_11_5  (
            .in0(N__19142),
            .in1(N__20491),
            .in2(N__19413),
            .in3(N__21564),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_6_o3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_9_11_6 .LUT_INIT=16'b1111010110100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_3_LC_9_11_6  (
            .in0(N__21071),
            .in1(N__23196),
            .in2(N__18902),
            .in3(N__20410),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_9_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_9_11_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_1_LC_9_11_7  (
            .in0(N__21365),
            .in1(_gnd_net_),
            .in2(N__18899),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.g1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_2_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_2_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_2_LC_9_12_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_2_LC_9_12_0  (
            .in0(N__23077),
            .in1(N__22862),
            .in2(_gnd_net_),
            .in3(N__22449),
            .lcout(\Lab_UT.dictrl.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_17_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_17_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_17_LC_9_12_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_17_LC_9_12_1  (
            .in0(N__20650),
            .in1(N__19064),
            .in2(N__21433),
            .in3(N__19049),
            .lcout(\Lab_UT.dictrl.N_16_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_5_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_5_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_5_LC_9_12_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_5_LC_9_12_2  (
            .in0(N__22556),
            .in1(N__22863),
            .in2(N__21571),
            .in3(N__22451),
            .lcout(\Lab_UT.dictrl.g0_i_a3_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_0_0_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_0_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_0_0_LC_9_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_0_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__21208),
            .in2(_gnd_net_),
            .in3(N__22610),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_6_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_6_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_6_LC_9_12_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_6_LC_9_12_4  (
            .in0(N__20482),
            .in1(N__19365),
            .in2(N__19220),
            .in3(N__23078),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_a3_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_14_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_14_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_14_LC_9_12_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_14_LC_9_12_5  (
            .in0(N__19607),
            .in1(N__23096),
            .in2(N__19217),
            .in3(N__19214),
            .lcout(\Lab_UT.dictrl.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state32_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state32_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state32_LC_9_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state32_LC_9_12_6  (
            .in0(N__22973),
            .in1(N__19093),
            .in2(N__22615),
            .in3(N__21247),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_4_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_4_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_4_LC_9_12_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_4_LC_9_12_7  (
            .in0(N__22450),
            .in1(N__20481),
            .in2(N__22557),
            .in3(N__22609),
            .lcout(\Lab_UT.dictrl.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_9_13_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_LC_9_13_0  (
            .in0(N__21210),
            .in1(N__19160),
            .in2(_gnd_net_),
            .in3(N__19141),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_23_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_23_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_23_LC_9_13_1 .LUT_INIT=16'b0111010011111100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_23_LC_9_13_1  (
            .in0(N__19094),
            .in1(N__21133),
            .in2(N__19067),
            .in3(N__19613),
            .lcout(\Lab_UT.dictrl.N_13_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_2_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_2_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_2_LC_9_13_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_2_2_LC_9_13_2  (
            .in0(N__22864),
            .in1(N__23073),
            .in2(_gnd_net_),
            .in3(N__22459),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_20_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_20_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_20_LC_9_13_3 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_20_LC_9_13_3  (
            .in0(N__19619),
            .in1(N__21134),
            .in2(N__19058),
            .in3(N__19055),
            .lcout(\Lab_UT.dictrl.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state32_1_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state32_1_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state32_1_LC_9_13_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state32_1_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__19449),
            .in2(_gnd_net_),
            .in3(N__19245),
            .lcout(\Lab_UT.dictrl.next_state32Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_3_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_3_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_3_LC_9_13_5 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_2_3_LC_9_13_5  (
            .in0(N__20462),
            .in1(N__21534),
            .in2(N__22972),
            .in3(N__22527),
            .lcout(\Lab_UT.dictrl.g1_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_1_1_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_1_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_1_1_LC_9_13_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.g0_1_1_LC_9_13_6  (
            .in0(N__22976),
            .in1(N__19450),
            .in2(N__22616),
            .in3(N__19246),
            .lcout(\Lab_UT.dictrl.g0_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_4_LC_9_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_4_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_4_LC_9_13_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_4_LC_9_13_7  (
            .in0(N__20463),
            .in1(N__19326),
            .in2(N__23086),
            .in3(N__21535),
            .lcout(\Lab_UT.dictrl.g0_i_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_LC_9_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_2_LC_9_14_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_2_LC_9_14_0  (
            .in0(N__19486),
            .in1(N__19601),
            .in2(N__22611),
            .in3(N__19552),
            .lcout(\Lab_UT.dictrl.g1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19324),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_fast_2_LC_9_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_9_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_9_14_2  (
            .in0(N__19323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_2_rep2_LC_9_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep2_LC_9_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep2_LC_9_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep2_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19325),
            .lcout(bu_rx_data_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_2_LC_9_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_9_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_14_4  (
            .in0(N__19322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19778),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_1_rep2_LC_9_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep2_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep2_LC_9_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_rep2_LC_9_14_7  (
            .in0(N__19779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22284),
            .ce(N__22074),
            .sr(N__22010));
    defparam \buart.Z_rx.shifter_3_rep1_LC_9_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_9_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22456),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22279),
            .ce(N__22072),
            .sr(N__22012));
    defparam \buart.Z_rx.shifter_fast_0_LC_9_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_9_15_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__22748),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22279),
            .ce(N__22072),
            .sr(N__22012));
    defparam \uu2.bitmap_34_LC_11_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_11_4_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_34_LC_11_4_4  (
            .in0(N__20066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20363),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__21953));
    defparam \uu2.bitmap_162_LC_11_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_11_4_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_162_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(N__19628),
            .in2(_gnd_net_),
            .in3(N__20065),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_34C_net ),
            .ce(),
            .sr(N__21953));
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_11_6_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_11_6_0 .LUT_INIT=16'b0111111101100111;
    LogicCell40 \Lab_UT.bcd2segment4.segment_0_2_LC_11_6_0  (
            .in0(N__20338),
            .in1(N__20272),
            .in2(N__20216),
            .in3(N__20144),
            .lcout(\Lab_UT.bcd2segment4.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_4_LC_11_6_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_4_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_4_LC_11_6_1 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_4_LC_11_6_1  (
            .in0(N__20213),
            .in1(N__20141),
            .in2(N__20274),
            .in3(N__20341),
            .lcout(\Lab_UT.bcd2segment4.segmentUQ_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_5_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_5_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_5_LC_11_6_2 .LUT_INIT=16'b1111100111011000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_5_LC_11_6_2  (
            .in0(N__20339),
            .in1(N__20264),
            .in2(N__20217),
            .in3(N__20145),
            .lcout(\Lab_UT.bcd2segment4.segmentUQ_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_6_LC_11_6_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_6_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_6_LC_11_6_3 .LUT_INIT=16'b1111100010100101;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_6_LC_11_6_3  (
            .in0(N__20214),
            .in1(N__20142),
            .in2(N__20275),
            .in3(N__20342),
            .lcout(\Lab_UT.bcd2segment4.segmentUQ_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_0_0_LC_11_6_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_0_0_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_0_0_LC_11_6_4 .LUT_INIT=16'b1011011011111101;
    LogicCell40 \Lab_UT.bcd2segment4.segment_0_0_LC_11_6_4  (
            .in0(N__20340),
            .in1(N__20268),
            .in2(N__20218),
            .in3(N__20146),
            .lcout(\Lab_UT.bcd2segment4.segment_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_11_6_5 .LUT_INIT=16'b0100100101111111;
    LogicCell40 \Lab_UT.bcd2segment4.segment_0_1_LC_11_6_5  (
            .in0(N__20215),
            .in1(N__20143),
            .in2(N__20276),
            .in3(N__20343),
            .lcout(\Lab_UT.bcd2segment4.segment_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_3_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_3_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_3_LC_11_6_6 .LUT_INIT=16'b1110110111001010;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_3_LC_11_6_6  (
            .in0(N__20344),
            .in1(N__20273),
            .in2(N__20219),
            .in3(N__20147),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_290_LC_11_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_11_6_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_290_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20069),
            .in3(N__20059),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__21951));
    defparam \Lab_UT.dictrl.state_0_3_rep1_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_LC_11_9_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_LC_11_9_0  (
            .in0(N__19908),
            .in1(N__20681),
            .in2(N__20866),
            .in3(N__21774),
            .lcout(\Lab_UT.dictrl.state_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__21988));
    defparam \Lab_UT.dictrl.state_0_fast_3_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_3_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_3_LC_11_9_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_3_LC_11_9_1  (
            .in0(N__21773),
            .in1(N__20865),
            .in2(N__20690),
            .in3(N__19910),
            .lcout(\Lab_UT.dictrl.state_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__21988));
    defparam \Lab_UT.dictrl.state_0_3_rep2_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_LC_11_9_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_LC_11_9_2  (
            .in0(N__19909),
            .in1(N__20682),
            .in2(N__20867),
            .in3(N__21775),
            .lcout(\Lab_UT.dictrl.state_3_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__21988));
    defparam \Lab_UT.dictrl.state_0_3_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_LC_11_9_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_LC_11_9_3  (
            .in0(N__21772),
            .in1(N__20858),
            .in2(N__20689),
            .in3(N__19907),
            .lcout(\Lab_UT.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22329),
            .ce(),
            .sr(N__21988));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_9_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_9_4  (
            .in0(N__20855),
            .in1(N__20601),
            .in2(N__21790),
            .in3(N__22036),
            .lcout(\Lab_UT.dictrl.g0_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_RNO_1_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_RNO_1_LC_11_9_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_RNO_1_LC_11_9_6  (
            .in0(N__20856),
            .in1(_gnd_net_),
            .in2(N__21791),
            .in3(N__20603),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_RNO_1_LC_11_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_1_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_RNO_1_LC_11_9_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_RNO_1_LC_11_9_7  (
            .in0(N__20602),
            .in1(N__20857),
            .in2(_gnd_net_),
            .in3(N__21768),
            .lcout(\Lab_UT.dictrl.g0_0_i_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_11_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_11_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m35_LC_11_10_7  (
            .in0(N__20732),
            .in1(N__20604),
            .in2(_gnd_net_),
            .in3(N__21605),
            .lcout(\Lab_UT.dictrl.N_40_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m12_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m12_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m12_LC_11_11_0 .LUT_INIT=16'b0010011100100010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m12_LC_11_11_0  (
            .in0(N__21130),
            .in1(N__20954),
            .in2(N__20662),
            .in3(N__21603),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m15_ns_LC_11_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m15_ns_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m15_ns_LC_11_11_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m15_ns_LC_11_11_1  (
            .in0(N__21455),
            .in1(_gnd_net_),
            .in2(N__20537),
            .in3(N__20420),
            .lcout(\Lab_UT.dictrl.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_6_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_6_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_6_LC_11_11_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_6_LC_11_11_2  (
            .in0(N__20512),
            .in1(N__20492),
            .in2(N__23087),
            .in3(N__21113),
            .lcout(\Lab_UT.dictrl.g1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_3_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_3_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_3_LC_11_11_3 .LUT_INIT=16'b0001001100010000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_3_LC_11_11_3  (
            .in0(N__21604),
            .in1(N__23170),
            .in2(N__21132),
            .in3(N__20409),
            .lcout(\Lab_UT.dictrl.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m20_LC_11_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m20_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m20_LC_11_11_4 .LUT_INIT=16'b0000011101010111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m20_LC_11_11_4  (
            .in0(N__21129),
            .in1(N__20408),
            .in2(N__23197),
            .in3(N__20953),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIFHHU6_2_LC_11_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIFHHU6_2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIFHHU6_2_LC_11_11_5 .LUT_INIT=16'b0001001110011011;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIFHHU6_2_LC_11_11_5  (
            .in0(N__21454),
            .in1(N__21764),
            .in2(N__21623),
            .in3(N__21280),
            .lcout(\Lab_UT.dictrl.next_state_latmux_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_11_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_11_11_6 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_11_11_6  (
            .in0(N__21182),
            .in1(N__21114),
            .in2(_gnd_net_),
            .in3(N__21602),
            .lcout(\Lab_UT.dictrl.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_LC_11_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_LC_11_11_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_1_LC_11_11_7  (
            .in0(N__22961),
            .in1(N__21568),
            .in2(N__22871),
            .in3(N__23083),
            .lcout(\Lab_UT.dictrl.g1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_11_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_11_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_11_12_0  (
            .in0(N__20909),
            .in1(N__21434),
            .in2(_gnd_net_),
            .in3(N__21281),
            .lcout(\Lab_UT.dictrl.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_11_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_11_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_1_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__23084),
            .in2(_gnd_net_),
            .in3(N__22434),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_LC_11_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_LC_11_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m17_LC_11_12_2  (
            .in0(N__22825),
            .in1(N__21140),
            .in2(N__21257),
            .in3(N__21254),
            .lcout(\Lab_UT.dictrl.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_1_LC_11_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m17_1_LC_11_12_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m17_1_LC_11_12_3  (
            .in0(N__22959),
            .in1(N__22599),
            .in2(N__21198),
            .in3(N__22502),
            .lcout(\Lab_UT.dictrl.m17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_5_LC_11_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_5_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_5_LC_11_12_4 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_5_LC_11_12_4  (
            .in0(N__23174),
            .in1(N__21131),
            .in2(_gnd_net_),
            .in3(N__20949),
            .lcout(\Lab_UT.dictrl.N_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_5_LC_11_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_5_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_5_LC_11_12_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_5_LC_11_12_5  (
            .in0(N__22960),
            .in1(N__22824),
            .in2(N__20899),
            .in3(N__22503),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_0_LC_11_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_0_LC_11_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_0_LC_11_12_6  (
            .in0(N__22435),
            .in1(N__22764),
            .in2(N__23231),
            .in3(N__23228),
            .lcout(\Lab_UT.dictrl.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_3_LC_11_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_3_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_3_LC_11_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_3_LC_11_12_7  (
            .in0(N__22826),
            .in1(N__22436),
            .in2(N__23198),
            .in3(N__22504),
            .lcout(\Lab_UT.dictrl.g0_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_11_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_11_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_6_LC_11_13_0  (
            .in0(N__23085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__22076),
            .sr(N__22011));
    defparam \buart.Z_rx.shifter_3_rep2_LC_11_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep2_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22419),
            .lcout(bu_rx_data_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__22076),
            .sr(N__22011));
    defparam \buart.Z_rx.shifter_5_LC_11_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22827),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22296),
            .ce(N__22076),
            .sr(N__22011));
    defparam \buart.Z_rx.shifter_0_rep1_LC_11_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_rep1_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22769),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22290),
            .ce(N__22075),
            .sr(N__22013));
    defparam \buart.Z_rx.shifter_4_LC_11_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22520),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22290),
            .ce(N__22075),
            .sr(N__22013));
endmodule // latticehx1k
