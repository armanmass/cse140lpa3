-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 20 2019 23:49:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu2.mem0.N_137\ : std_logic;
signal \uu2.mem0.N_141\ : std_logic;
signal \uu2.bitmap_pmux_u_0_a2_0_cascade_\ : std_logic;
signal \uu2.mem0.N_140\ : std_logic;
signal \uu2.mem0.N_139\ : std_logic;
signal \INVuu2.w_addr_user_1C_net\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.un4_l_count_16_cascade_\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un55_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_0_8_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu2.N_34_cascade_\ : std_logic;
signal \uu2.N_114\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.mem0.N_31_i\ : std_logic;
signal \uu2.mem0.N_61_cascade_\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.N_922_tz_tz\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \uu2.bitmap_pmux_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.N_37\ : std_logic;
signal \uu2.mem0.N_59\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.un404_ci_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \INVuu2.w_addr_user_4C_net\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu2.un1_l_count_2_2_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.un306_ci_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu2.w_data_0_a2_0_6_cascade_\ : std_logic;
signal \uu2.w_data_0_a2_2_6\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_4C_net\ : std_logic;
signal \uu2.bitmap_pmux_u_0_a2_0_2_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_2C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \INVuu2.bitmap_186C_net\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmap_RNIRETJ1Z0Z_93_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1_cascade_\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \uu2.mem0.N_135\ : std_logic;
signal \uu2.mem0.N_134\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_7C_net\ : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_\ : std_logic;
signal \uu2.N_32_0\ : std_logic;
signal \uu2.mem0.N_133\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.N_161_cascade_\ : std_logic;
signal \INVuu2.w_addr_user_nesr_8C_net\ : std_logic;
signal \uu2.N_101_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.N_106_cascade_\ : std_logic;
signal \uu2.N_164\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_3_6\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_2_6_cascade_\ : std_logic;
signal \uu2.N_230\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.mem0.N_138\ : std_logic;
signal \oneSecStrb_cascade_\ : std_logic;
signal clk : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.N_102\ : std_logic;
signal \uu2.mem0.N_54_i\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.bitmap_pmux_25_i_m2_am_1_cascade_\ : std_logic;
signal \uu2.bitmap_RNIG91I1Z0Z_66\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \INVuu2.bitmap_194C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.N_34\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.N_47\ : std_logic;
signal \uu2.N_38\ : std_logic;
signal \uu2.w_addr_displaying_RNI0ES07Z0Z_5\ : std_logic;
signal \uu2.N_33\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_3_rep1C_net\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.mem0.N_136\ : std_logic;
signal \uu2.bitmap_RNIFJI02Z0Z_212\ : std_logic;
signal \uu2.N_65\ : std_logic;
signal \uu2.bitmap_pmux_u_0_83_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.N_112_i\ : std_logic;
signal \uu2.N_100_cascade_\ : std_logic;
signal \uu2.N_921_tz_tz\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.N_923_tz_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI8ND5GZ0Z_3\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmap_pmux_25_i_m2_bm_1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.bitmap_pmux_21_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.N_393_cascade_\ : std_logic;
signal \uu2.N_397\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.N_128\ : std_logic;
signal \uu2.N_131\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.sec2_1\ : std_logic;
signal \Lab_UT.sec2_2\ : std_logic;
signal \Lab_UT.sec2_3\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_a2_0Z0Z_4\ : std_logic;
signal \Lab_UT.dispString.un42_dOutP_cascade_\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_a2_0Z0Z_0\ : std_logic;
signal \Lab_UT.dispString.N_211_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_2\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \uu2.un1_w_user_cr_0\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_191\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3\ : std_logic;
signal \buart.Z_rx.idle_0_cascade_\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_rx.valid_1_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \INVuu2.bitmap_168C_net\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmap_pmux_24_bm_1\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.bitmap_RNI5T9T1Z0Z_72\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux\ : std_logic;
signal \uu2.N_237\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15\ : std_logic;
signal \uu2.N_395_cascade_\ : std_logic;
signal \uu2.N_401\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmap_pmux_15_i_m2_ns_1\ : std_logic;
signal \uu2.N_123\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.bitmap_RNIU2ISZ0Z_52\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.bitmap_pmux_24_am_1\ : std_logic;
signal \Lab_UT.min1_1\ : std_logic;
signal \Lab_UT.dispString.un46_dOutP_2\ : std_logic;
signal \Lab_UT.sec2_0\ : std_logic;
signal \G_190\ : std_logic;
signal \G_190_cascade_\ : std_logic;
signal \Lab_UT.dispString.i21_mux\ : std_logic;
signal \Lab_UT.dispString.m28_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_204\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.N_106\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \INVuu2.w_addr_user_nesr_5C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_0\ : std_logic;
signal \G_193\ : std_logic;
signal \G_193_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_219\ : std_logic;
signal \Lab_UT.dispString.N_222_cascade_\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \G_189\ : std_logic;
signal \G_189_cascade_\ : std_logic;
signal \Lab_UT.dispString.un42_dOutP\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \uu0_sec_clkD\ : std_logic;
signal \Lab_UT.dispString.m44_ns_1\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \Lab_UT.dispString.m42_ns_1\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \Lab_UT.dictrl.g1Z0Z_5\ : std_logic;
signal \Lab_UT.dictrl.g1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_2_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_1_7\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_1Z0Z_6\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_1_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_2\ : std_logic;
signal \Lab_UT.dictrl.N_19\ : std_logic;
signal \Lab_UT.dictrl.g0_17_o6_1Z0Z_5\ : std_logic;
signal \Lab_UT.min2_3\ : std_logic;
signal \Lab_UT.min1_3\ : std_logic;
signal \Lab_UT.min1_2\ : std_logic;
signal \Lab_UT.min1_0\ : std_logic;
signal \Lab_UT.min2_1\ : std_logic;
signal \Lab_UT.min2_0\ : std_logic;
signal \Lab_UT.min2_2\ : std_logic;
signal \Lab_UT.dispString.N_18_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_0Z0Z_1\ : std_logic;
signal \uu2.N_101\ : std_logic;
signal \uu2.N_111\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \Lab_UT.sec1_2\ : std_logic;
signal \Lab_UT.sec1_1\ : std_logic;
signal \Lab_UT.sec1_0\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \INVuu2.w_addr_user_7C_net\ : std_logic;
signal \Lab_UT.sec1_3\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_1\ : std_logic;
signal \Lab_UT.didp.countrce4.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_95_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_21_0_cascade_\ : std_logic;
signal \Lab_UT.i16_mux\ : std_logic;
signal \Lab_UT.dictrl.i18_mux\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_1Z0Z_1\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.dispString.m49_ns_1\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.un1_idle_1_0_iclkZ0\ : std_logic;
signal \G_186_cascade_\ : std_logic;
signal \G_191\ : std_logic;
signal \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_10_1\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dicRun_2\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_90_0\ : std_logic;
signal \Lab_UT.dictrl.N_95_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.LdStens_i_3\ : std_logic;
signal \Lab_UT.dictrl.state_fast_1\ : std_logic;
signal \Lab_UT.dictrl.N_95_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_5\ : std_logic;
signal \Lab_UT.dictrl.g0_2Z0Z_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0\ : std_logic;
signal \Lab_UT.dictrl.g1_1\ : std_logic;
signal \Lab_UT.dictrl.g2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_90_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.m40_N_5_mux_0\ : std_logic;
signal \Lab_UT.dictrl.g2Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_2_1\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_3_6\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_3_8\ : std_logic;
signal \Lab_UT.dictrl.N_22_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_17_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_0\ : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal \Lab_UT.didp.reset_12_1_3\ : std_logic;
signal \Lab_UT.didp.di_Mtens_2\ : std_logic;
signal \Lab_UT.didp.ce_12_3_cascade_\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.didp.un24_ce_2\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMtens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_1\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_0\ : std_logic;
signal \Lab_UT.didp.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.di_Stens_1\ : std_logic;
signal \Lab_UT.didp.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.regrce3.did_alarmMatch_3\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_0\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_1_cascade_\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_2\ : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_7\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_4_cascade_\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_5\ : std_logic;
signal \Lab_UT.did_alarmMatch_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_0_cascade_\ : std_logic;
signal \Lab_UT.did_alarmMatch_13\ : std_logic;
signal \G_183_cascade_\ : std_logic;
signal \Lab_UT.did_alarmMatch_12\ : std_logic;
signal \Lab_UT.didp.countrce2.un13_qPone\ : std_logic;
signal \Lab_UT.didp.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_2\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\ : std_logic;
signal \G_184\ : std_logic;
signal \Lab_UT.alarmstate_0_sqmuxa_1\ : std_logic;
signal \Lab_UT.didp.countrce1.un13_qPone\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.un1_armed_2_0_iso_iZ0\ : std_logic;
signal \Lab_UT.un1_idle_5_0_iclkZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.un1_armed_2_0_iso_iZ0_cascade_\ : std_logic;
signal \G_192\ : std_logic;
signal \Lab_UT.dictrl.N_113_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_fast_2\ : std_logic;
signal \Lab_UT.dictrl.g0_17_0\ : std_logic;
signal \Lab_UT.dictrl.g0_17_1\ : std_logic;
signal \Lab_UT.didp.di_Sones_2\ : std_logic;
signal \Lab_UT.didp.di_Sones_3\ : std_logic;
signal \Lab_UT.didp.un18_ce\ : std_logic;
signal \Lab_UT.LdSones_i_3\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.LdStens\ : std_logic;
signal bu_rx_data_rdy_0_g : std_logic;
signal \Lab_UT.dictrl.m30_0Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m25Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m59_ns_1_xZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.N_81_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_113_1\ : std_logic;
signal \Lab_UT.dictrl.N_113_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m59_ns_1\ : std_logic;
signal \Lab_UT.dictrl.N_81_0\ : std_logic;
signal \Lab_UT.dictrl.N_16_mux_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_113_0_0\ : std_logic;
signal \Lab_UT.dictrl.state_2_rep1\ : std_logic;
signal \Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5_0\ : std_logic;
signal \Lab_UT.dictrl.g2_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_0\ : std_logic;
signal \Lab_UT.dictrl.N_77_0\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep1\ : std_logic;
signal \Lab_UT.dictrl.g0_0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_2Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_77_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_77_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_2353_0_0\ : std_logic;
signal \buart__rx_shifter_fast_6\ : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \Lab_UT.dictrl.state_fast_3\ : std_logic;
signal \Lab_UT.dictrl.g1_6\ : std_logic;
signal \Lab_UT.dictrl.m47_xZ0Z0_cascade_\ : std_logic;
signal bu_rx_data_fast_4 : std_logic;
signal \Lab_UT.dictrl.m30Z0Z_1\ : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \Lab_UT.dictrl.g1_1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g2_1_0\ : std_logic;
signal \Lab_UT.dictrl.g2\ : std_logic;
signal \Lab_UT.didp.countrce3.ce_12_2_3\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.didp.regrce4.LdAMtens_0\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.didp.di_Mtens_0\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_6\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0\ : std_logic;
signal \Lab_UT.didp.di_Mones_3\ : std_logic;
signal \Lab_UT.didp.di_Mones_0\ : std_logic;
signal \Lab_UT.didp.di_Mones_1\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mones_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.N_13_0\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \G_183\ : std_logic;
signal \G_185\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m3_0\ : std_logic;
signal \Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_\ : std_logic;
signal \G_188\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8Z0Z_3\ : std_logic;
signal \G_188_cascade_\ : std_logic;
signal \G_187\ : std_logic;
signal \G_186\ : std_logic;
signal \G_187_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\ : std_logic;
signal \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\ : std_logic;
signal \Lab_UT.state_i_3_0\ : std_logic;
signal \Lab_UT.dictrl.g0_2Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m40_N_5_mux_1\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8Z0Z_4\ : std_logic;
signal \Lab_UT.didp.di_Sones_0\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal \Lab_UT.didp.di_Sones_1\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1\ : std_logic;
signal \Lab_UT.dictrl.N_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_12\ : std_logic;
signal \Lab_UT.dictrl.N_81\ : std_logic;
signal \Lab_UT.dictrl.next_state_i_1_2\ : std_logic;
signal \Lab_UT.dictrl.P8_mux\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_3\ : std_logic;
signal \Lab_UT.dictrl.P6_mux_0\ : std_logic;
signal \Lab_UT.dictrl.state_i_3_2\ : std_logic;
signal \Lab_UT.dictrl.N_114_mux\ : std_logic;
signal \Lab_UT.dictrl.N_69\ : std_logic;
signal \Lab_UT.dictrl.i10_mux\ : std_logic;
signal \Lab_UT.dictrl.N_69_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_0_3\ : std_logic;
signal \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_0_1\ : std_logic;
signal \Lab_UT.dictrl.P6_mux\ : std_logic;
signal \Lab_UT.dictrl.N_189\ : std_logic;
signal \Lab_UT.dictrl.m40_N_5_mux\ : std_logic;
signal \Lab_UT.dictrl.N_77\ : std_logic;
signal \Lab_UT.dictrl.N_77_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m73Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.m77_ns_1\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_106_mux\ : std_logic;
signal \Lab_UT.dictrl.m51_0\ : std_logic;
signal \Lab_UT.dictrl.state_i_3_1\ : std_logic;
signal \Lab_UT.dictrl.N_118_mux_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_3_1_1\ : std_logic;
signal \Lab_UT.dictrl.g0_17_a6_3Z0Z_7\ : std_logic;
signal \buart__rx_shifter_fast_0\ : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal \buart__rx_shifter_fast_5\ : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal \Lab_UT.dictrl.N_103_mux\ : std_logic;
signal \Lab_UT.dictrl.N_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_1_rep1\ : std_logic;
signal \Lab_UT.dictrl.N_12_0\ : std_logic;
signal \Lab_UT.LdASones\ : std_logic;
signal \Lab_UT.didp.regrce1.LdASones_0\ : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \shifter_7_rep1_RNIG7Q01\ : std_logic;
signal \buart.Z_rx.P7_mux\ : std_logic;
signal \N_16_mux\ : std_logic;
signal \shifter_7_rep1_RNIG7Q01_cascade_\ : std_logic;
signal \N_97\ : std_logic;
signal bu_rx_data_4_rep1 : std_logic;
signal bu_rx_data_rdy_0 : std_logic;
signal \Lab_UT_dictrl_state_3_rep2\ : std_logic;
signal \Lab_UT.dictrl.g0_5_a4_1_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_90\ : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal rst_g : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.dictrl.m25Z0Z_0\ : std_logic;
signal \N_119_mux_cascade_\ : std_logic;
signal bu_rx_data_3_rep2 : std_logic;
signal \Lab_UT.dictrl.g0_5_a4_1_4\ : std_logic;
signal \Lab_UT.dictrl.m86Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m86Z0Z_2\ : std_logic;
signal \Lab_UT.state_3\ : std_logic;
signal \Lab_UT.dictrl.un1_next_state66_0\ : std_logic;
signal \Lab_UT.state_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_1_a0_0_0\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_4 : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.dictrl.g0_5_o4_3\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.g0_5_o4_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_11\ : std_logic;
signal \N_117_cascade_\ : std_logic;
signal \resetGen_reset_count_0\ : std_logic;
signal \resetGen_reset_count_1\ : std_logic;
signal \resetGen_reset_count_2_2_cascade_\ : std_logic;
signal \resetGen_reset_count_2\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \N_91_i\ : std_logic;
signal clk_g : std_logic;
signal \N_119_mux\ : std_logic;
signal \resetGen_reset_count_4\ : std_logic;
signal m87 : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__8436\&\N__8412\&\N__8385\&\N__8475\&\N__8538\&\N__8361\&\N__8328\&\N__8577\&\N__8619\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__9489\&\N__9528\&\N__9540\&\N__10239\&\N__7725\&\N__9777\&\N__7752\&\N__7698\&\N__7713\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__8103\&'0'&\N__8295\&'0'&\N__8280\&'0'&\N__8259\&'0'&\N__9981\&'0'&\N__8286\&'0'&\N__8229\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__7686\,
            RESETB => \N__15729\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21667\,
            RE => \N__15744\,
            WCLKE => \N__9737\,
            WCLK => \N__21666\,
            WE => \N__9738\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21862\,
            DIN => \N__21861\,
            DOUT => \N__21860\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__21862\,
            PADOUT => \N__21861\,
            PADIN => \N__21860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21853\,
            DIN => \N__21852\,
            DOUT => \N__21851\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__21853\,
            PADOUT => \N__21852\,
            PADIN => \N__21851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21844\,
            DIN => \N__21843\,
            DOUT => \N__21842\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__21844\,
            PADOUT => \N__21843\,
            PADIN => \N__21842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21835\,
            DIN => \N__21834\,
            DOUT => \N__21833\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21835\,
            PADOUT => \N__21834\,
            PADIN => \N__21833\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__21630\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21826\,
            DIN => \N__21825\,
            DOUT => \N__21824\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21826\,
            PADOUT => \N__21825\,
            PADIN => \N__21824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21817\,
            DIN => \N__21816\,
            DOUT => \N__21815\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__21817\,
            PADOUT => \N__21816\,
            PADIN => \N__21815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21808\,
            DIN => \N__21807\,
            DOUT => \N__21806\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__21808\,
            PADOUT => \N__21807\,
            PADIN => \N__21806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21799\,
            DIN => \N__21798\,
            DOUT => \N__21797\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21799\,
            PADOUT => \N__21798\,
            PADIN => \N__21797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21790\,
            DIN => \N__21789\,
            DOUT => \N__21788\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21790\,
            PADOUT => \N__21789\,
            PADIN => \N__21788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21781\,
            DIN => \N__21780\,
            DOUT => \N__21779\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21781\,
            PADOUT => \N__21780\,
            PADIN => \N__21779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__21762\,
            I => \N_117_cascade_\
        );

    \I__5344\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21752\
        );

    \I__5343\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21743\
        );

    \I__5342\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21743\
        );

    \I__5341\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21743\
        );

    \I__5340\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21743\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__21752\,
            I => \resetGen_reset_count_0\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__21743\,
            I => \resetGen_reset_count_0\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__21738\,
            I => \N__21734\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__21737\,
            I => \N__21731\
        );

    \I__5335\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21720\
        );

    \I__5334\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21720\
        );

    \I__5333\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21720\
        );

    \I__5332\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21720\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__21720\,
            I => \resetGen_reset_count_1\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__21717\,
            I => \resetGen_reset_count_2_2_cascade_\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__21714\,
            I => \N__21708\
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__21713\,
            I => \N__21705\
        );

    \I__5327\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21696\
        );

    \I__5326\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21696\
        );

    \I__5325\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21696\
        );

    \I__5324\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21696\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__21696\,
            I => \resetGen_reset_count_2\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__5321\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21684\
        );

    \I__5320\ : InMux
    port map (
            O => \N__21689\,
            I => \N__21684\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__21684\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__5318\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21675\
        );

    \I__5317\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21675\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__21675\,
            I => \N_91_i\
        );

    \I__5315\ : ClkMux
    port map (
            O => \N__21672\,
            I => \N__21429\
        );

    \I__5314\ : ClkMux
    port map (
            O => \N__21671\,
            I => \N__21429\
        );

    \I__5313\ : ClkMux
    port map (
            O => \N__21670\,
            I => \N__21429\
        );

    \I__5312\ : ClkMux
    port map (
            O => \N__21669\,
            I => \N__21429\
        );

    \I__5311\ : ClkMux
    port map (
            O => \N__21668\,
            I => \N__21429\
        );

    \I__5310\ : ClkMux
    port map (
            O => \N__21667\,
            I => \N__21429\
        );

    \I__5309\ : ClkMux
    port map (
            O => \N__21666\,
            I => \N__21429\
        );

    \I__5308\ : ClkMux
    port map (
            O => \N__21665\,
            I => \N__21429\
        );

    \I__5307\ : ClkMux
    port map (
            O => \N__21664\,
            I => \N__21429\
        );

    \I__5306\ : ClkMux
    port map (
            O => \N__21663\,
            I => \N__21429\
        );

    \I__5305\ : ClkMux
    port map (
            O => \N__21662\,
            I => \N__21429\
        );

    \I__5304\ : ClkMux
    port map (
            O => \N__21661\,
            I => \N__21429\
        );

    \I__5303\ : ClkMux
    port map (
            O => \N__21660\,
            I => \N__21429\
        );

    \I__5302\ : ClkMux
    port map (
            O => \N__21659\,
            I => \N__21429\
        );

    \I__5301\ : ClkMux
    port map (
            O => \N__21658\,
            I => \N__21429\
        );

    \I__5300\ : ClkMux
    port map (
            O => \N__21657\,
            I => \N__21429\
        );

    \I__5299\ : ClkMux
    port map (
            O => \N__21656\,
            I => \N__21429\
        );

    \I__5298\ : ClkMux
    port map (
            O => \N__21655\,
            I => \N__21429\
        );

    \I__5297\ : ClkMux
    port map (
            O => \N__21654\,
            I => \N__21429\
        );

    \I__5296\ : ClkMux
    port map (
            O => \N__21653\,
            I => \N__21429\
        );

    \I__5295\ : ClkMux
    port map (
            O => \N__21652\,
            I => \N__21429\
        );

    \I__5294\ : ClkMux
    port map (
            O => \N__21651\,
            I => \N__21429\
        );

    \I__5293\ : ClkMux
    port map (
            O => \N__21650\,
            I => \N__21429\
        );

    \I__5292\ : ClkMux
    port map (
            O => \N__21649\,
            I => \N__21429\
        );

    \I__5291\ : ClkMux
    port map (
            O => \N__21648\,
            I => \N__21429\
        );

    \I__5290\ : ClkMux
    port map (
            O => \N__21647\,
            I => \N__21429\
        );

    \I__5289\ : ClkMux
    port map (
            O => \N__21646\,
            I => \N__21429\
        );

    \I__5288\ : ClkMux
    port map (
            O => \N__21645\,
            I => \N__21429\
        );

    \I__5287\ : ClkMux
    port map (
            O => \N__21644\,
            I => \N__21429\
        );

    \I__5286\ : ClkMux
    port map (
            O => \N__21643\,
            I => \N__21429\
        );

    \I__5285\ : ClkMux
    port map (
            O => \N__21642\,
            I => \N__21429\
        );

    \I__5284\ : ClkMux
    port map (
            O => \N__21641\,
            I => \N__21429\
        );

    \I__5283\ : ClkMux
    port map (
            O => \N__21640\,
            I => \N__21429\
        );

    \I__5282\ : ClkMux
    port map (
            O => \N__21639\,
            I => \N__21429\
        );

    \I__5281\ : ClkMux
    port map (
            O => \N__21638\,
            I => \N__21429\
        );

    \I__5280\ : ClkMux
    port map (
            O => \N__21637\,
            I => \N__21429\
        );

    \I__5279\ : ClkMux
    port map (
            O => \N__21636\,
            I => \N__21429\
        );

    \I__5278\ : ClkMux
    port map (
            O => \N__21635\,
            I => \N__21429\
        );

    \I__5277\ : ClkMux
    port map (
            O => \N__21634\,
            I => \N__21429\
        );

    \I__5276\ : ClkMux
    port map (
            O => \N__21633\,
            I => \N__21429\
        );

    \I__5275\ : ClkMux
    port map (
            O => \N__21632\,
            I => \N__21429\
        );

    \I__5274\ : ClkMux
    port map (
            O => \N__21631\,
            I => \N__21429\
        );

    \I__5273\ : ClkMux
    port map (
            O => \N__21630\,
            I => \N__21429\
        );

    \I__5272\ : ClkMux
    port map (
            O => \N__21629\,
            I => \N__21429\
        );

    \I__5271\ : ClkMux
    port map (
            O => \N__21628\,
            I => \N__21429\
        );

    \I__5270\ : ClkMux
    port map (
            O => \N__21627\,
            I => \N__21429\
        );

    \I__5269\ : ClkMux
    port map (
            O => \N__21626\,
            I => \N__21429\
        );

    \I__5268\ : ClkMux
    port map (
            O => \N__21625\,
            I => \N__21429\
        );

    \I__5267\ : ClkMux
    port map (
            O => \N__21624\,
            I => \N__21429\
        );

    \I__5266\ : ClkMux
    port map (
            O => \N__21623\,
            I => \N__21429\
        );

    \I__5265\ : ClkMux
    port map (
            O => \N__21622\,
            I => \N__21429\
        );

    \I__5264\ : ClkMux
    port map (
            O => \N__21621\,
            I => \N__21429\
        );

    \I__5263\ : ClkMux
    port map (
            O => \N__21620\,
            I => \N__21429\
        );

    \I__5262\ : ClkMux
    port map (
            O => \N__21619\,
            I => \N__21429\
        );

    \I__5261\ : ClkMux
    port map (
            O => \N__21618\,
            I => \N__21429\
        );

    \I__5260\ : ClkMux
    port map (
            O => \N__21617\,
            I => \N__21429\
        );

    \I__5259\ : ClkMux
    port map (
            O => \N__21616\,
            I => \N__21429\
        );

    \I__5258\ : ClkMux
    port map (
            O => \N__21615\,
            I => \N__21429\
        );

    \I__5257\ : ClkMux
    port map (
            O => \N__21614\,
            I => \N__21429\
        );

    \I__5256\ : ClkMux
    port map (
            O => \N__21613\,
            I => \N__21429\
        );

    \I__5255\ : ClkMux
    port map (
            O => \N__21612\,
            I => \N__21429\
        );

    \I__5254\ : ClkMux
    port map (
            O => \N__21611\,
            I => \N__21429\
        );

    \I__5253\ : ClkMux
    port map (
            O => \N__21610\,
            I => \N__21429\
        );

    \I__5252\ : ClkMux
    port map (
            O => \N__21609\,
            I => \N__21429\
        );

    \I__5251\ : ClkMux
    port map (
            O => \N__21608\,
            I => \N__21429\
        );

    \I__5250\ : ClkMux
    port map (
            O => \N__21607\,
            I => \N__21429\
        );

    \I__5249\ : ClkMux
    port map (
            O => \N__21606\,
            I => \N__21429\
        );

    \I__5248\ : ClkMux
    port map (
            O => \N__21605\,
            I => \N__21429\
        );

    \I__5247\ : ClkMux
    port map (
            O => \N__21604\,
            I => \N__21429\
        );

    \I__5246\ : ClkMux
    port map (
            O => \N__21603\,
            I => \N__21429\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__21602\,
            I => \N__21429\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__21601\,
            I => \N__21429\
        );

    \I__5243\ : ClkMux
    port map (
            O => \N__21600\,
            I => \N__21429\
        );

    \I__5242\ : ClkMux
    port map (
            O => \N__21599\,
            I => \N__21429\
        );

    \I__5241\ : ClkMux
    port map (
            O => \N__21598\,
            I => \N__21429\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__21597\,
            I => \N__21429\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__21596\,
            I => \N__21429\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__21595\,
            I => \N__21429\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__21594\,
            I => \N__21429\
        );

    \I__5236\ : ClkMux
    port map (
            O => \N__21593\,
            I => \N__21429\
        );

    \I__5235\ : ClkMux
    port map (
            O => \N__21592\,
            I => \N__21429\
        );

    \I__5234\ : GlobalMux
    port map (
            O => \N__21429\,
            I => \N__21426\
        );

    \I__5233\ : gio2CtrlBuf
    port map (
            O => \N__21426\,
            I => clk_g
        );

    \I__5232\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21402\
        );

    \I__5231\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21402\
        );

    \I__5230\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21402\
        );

    \I__5229\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21402\
        );

    \I__5228\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21402\
        );

    \I__5227\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21402\
        );

    \I__5226\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21402\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N_119_mux\
        );

    \I__5224\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21393\
        );

    \I__5223\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21388\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21383\
        );

    \I__5221\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21383\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__21393\,
            I => \N__21380\
        );

    \I__5219\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21375\
        );

    \I__5218\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21375\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__21388\,
            I => \resetGen_reset_count_4\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__21383\,
            I => \resetGen_reset_count_4\
        );

    \I__5215\ : Odrv12
    port map (
            O => \N__21380\,
            I => \resetGen_reset_count_4\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__21375\,
            I => \resetGen_reset_count_4\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__21363\,
            I => m87
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__21360\,
            I => \N_119_mux_cascade_\
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__21357\,
            I => \N__21352\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__21356\,
            I => \N__21349\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__21355\,
            I => \N__21345\
        );

    \I__5207\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21342\
        );

    \I__5206\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21339\
        );

    \I__5205\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21334\
        );

    \I__5204\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21334\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__21342\,
            I => \N__21329\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__21339\,
            I => \N__21321\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__21334\,
            I => \N__21318\
        );

    \I__5200\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21313\
        );

    \I__5199\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21313\
        );

    \I__5198\ : Span4Mux_s2_h
    port map (
            O => \N__21329\,
            I => \N__21310\
        );

    \I__5197\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21305\
        );

    \I__5196\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21305\
        );

    \I__5195\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21302\
        );

    \I__5194\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21297\
        );

    \I__5193\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21297\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__21321\,
            I => \N__21292\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__21318\,
            I => \N__21292\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21289\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__21310\,
            I => bu_rx_data_3_rep2
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__21305\,
            I => bu_rx_data_3_rep2
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__21302\,
            I => bu_rx_data_3_rep2
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__21297\,
            I => bu_rx_data_3_rep2
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__21292\,
            I => bu_rx_data_3_rep2
        );

    \I__5184\ : Odrv12
    port map (
            O => \N__21289\,
            I => bu_rx_data_3_rep2
        );

    \I__5183\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__21273\,
            I => \Lab_UT.dictrl.g0_5_a4_1_4\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__21270\,
            I => \Lab_UT.dictrl.m86Z0Z_0_cascade_\
        );

    \I__5180\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21264\,
            I => \Lab_UT.dictrl.m86Z0Z_2\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__21261\,
            I => \N__21256\
        );

    \I__5177\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21252\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__21259\,
            I => \N__21247\
        );

    \I__5175\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21244\
        );

    \I__5174\ : CascadeMux
    port map (
            O => \N__21255\,
            I => \N__21240\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21233\
        );

    \I__5172\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21230\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21227\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21224\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21221\
        );

    \I__5168\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21218\
        );

    \I__5167\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21213\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__21239\,
            I => \N__21208\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__21238\,
            I => \N__21205\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__21237\,
            I => \N__21201\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21198\
        );

    \I__5162\ : Span4Mux_v
    port map (
            O => \N__21233\,
            I => \N__21191\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__21230\,
            I => \N__21191\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__21227\,
            I => \N__21188\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21185\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__21221\,
            I => \N__21180\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21180\
        );

    \I__5156\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21177\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__21216\,
            I => \N__21173\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__21213\,
            I => \N__21170\
        );

    \I__5153\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21165\
        );

    \I__5152\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21165\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21160\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21160\
        );

    \I__5149\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21155\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21155\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__21198\,
            I => \N__21152\
        );

    \I__5146\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21149\
        );

    \I__5145\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21146\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__21191\,
            I => \N__21141\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__21188\,
            I => \N__21141\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__21185\,
            I => \N__21134\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__21180\,
            I => \N__21134\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21134\
        );

    \I__5139\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21129\
        );

    \I__5138\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21129\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__21170\,
            I => \N__21122\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__21165\,
            I => \N__21122\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21122\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21155\,
            I => \Lab_UT.state_3\
        );

    \I__5133\ : Odrv12
    port map (
            O => \N__21152\,
            I => \Lab_UT.state_3\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__21149\,
            I => \Lab_UT.state_3\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__21146\,
            I => \Lab_UT.state_3\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__21141\,
            I => \Lab_UT.state_3\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__21134\,
            I => \Lab_UT.state_3\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__21129\,
            I => \Lab_UT.state_3\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__21122\,
            I => \Lab_UT.state_3\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21093\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__21104\,
            I => \N__21088\
        );

    \I__5124\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21085\
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__21102\,
            I => \N__21080\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21075\
        );

    \I__5121\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21072\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21065\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21065\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21065\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21062\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21093\,
            I => \N__21059\
        );

    \I__5115\ : CascadeMux
    port map (
            O => \N__21092\,
            I => \N__21053\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__21091\,
            I => \N__21050\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21045\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21041\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21032\
        );

    \I__5110\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21032\
        );

    \I__5109\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21032\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21032\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21029\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21075\,
            I => \N__21024\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21024\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__21065\,
            I => \N__21013\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21062\,
            I => \N__21013\
        );

    \I__5102\ : Span4Mux_s1_h
    port map (
            O => \N__21059\,
            I => \N__21013\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21002\
        );

    \I__5100\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21002\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21002\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21002\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21002\
        );

    \I__5096\ : InMux
    port map (
            O => \N__21049\,
            I => \N__20997\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21048\,
            I => \N__20997\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__21045\,
            I => \N__20994\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__21044\,
            I => \N__20991\
        );

    \I__5092\ : Span4Mux_v
    port map (
            O => \N__21041\,
            I => \N__20988\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__20981\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__20981\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__21024\,
            I => \N__20981\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21023\,
            I => \N__20978\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21022\,
            I => \N__20975\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21021\,
            I => \N__20970\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21020\,
            I => \N__20970\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__21013\,
            I => \N__20967\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20964\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__20997\,
            I => \N__20959\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__20994\,
            I => \N__20959\
        );

    \I__5080\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20956\
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__20988\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__20981\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__20978\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__20975\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__20970\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__20967\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__20964\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__20959\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__20956\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__20937\,
            I => \N__20931\
        );

    \I__5069\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20920\
        );

    \I__5068\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20917\
        );

    \I__5067\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20914\
        );

    \I__5066\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20911\
        );

    \I__5065\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20908\
        );

    \I__5064\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20903\
        );

    \I__5063\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20894\
        );

    \I__5062\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20894\
        );

    \I__5061\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20894\
        );

    \I__5060\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20894\
        );

    \I__5059\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20888\
        );

    \I__5058\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20888\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20874\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20871\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20866\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__20911\,
            I => \N__20866\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20863\
        );

    \I__5052\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20858\
        );

    \I__5051\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20858\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20855\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20852\
        );

    \I__5048\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20849\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20846\
        );

    \I__5046\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20843\
        );

    \I__5045\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20840\
        );

    \I__5044\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20831\
        );

    \I__5043\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20831\
        );

    \I__5042\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20831\
        );

    \I__5041\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20831\
        );

    \I__5040\ : InMux
    port map (
            O => \N__20881\,
            I => \N__20828\
        );

    \I__5039\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20823\
        );

    \I__5038\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20823\
        );

    \I__5037\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20818\
        );

    \I__5036\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20818\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__20874\,
            I => \N__20815\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__20871\,
            I => \N__20810\
        );

    \I__5033\ : Span4Mux_v
    port map (
            O => \N__20866\,
            I => \N__20810\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__20863\,
            I => \N__20803\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__20858\,
            I => \N__20803\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__20855\,
            I => \N__20803\
        );

    \I__5029\ : Span4Mux_s3_h
    port map (
            O => \N__20852\,
            I => \N__20796\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__20849\,
            I => \N__20796\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__20846\,
            I => \N__20796\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__20843\,
            I => \Lab_UT.state_0\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__20840\,
            I => \Lab_UT.state_0\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__20831\,
            I => \Lab_UT.state_0\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__20828\,
            I => \Lab_UT.state_0\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__20823\,
            I => \Lab_UT.state_0\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__20818\,
            I => \Lab_UT.state_0\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__20815\,
            I => \Lab_UT.state_0\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__20810\,
            I => \Lab_UT.state_0\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__20803\,
            I => \Lab_UT.state_0\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__20796\,
            I => \Lab_UT.state_0\
        );

    \I__5016\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__5014\ : Odrv12
    port map (
            O => \N__20769\,
            I => \Lab_UT.dictrl.next_state_latmux_1_a0_0_0\
        );

    \I__5013\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20761\
        );

    \I__5012\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20758\
        );

    \I__5011\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20749\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20744\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20744\
        );

    \I__5008\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20734\
        );

    \I__5007\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20734\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \N__20728\
        );

    \I__5005\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20725\
        );

    \I__5004\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20722\
        );

    \I__5003\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20719\
        );

    \I__5002\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20716\
        );

    \I__5001\ : Span4Mux_v
    port map (
            O => \N__20744\,
            I => \N__20713\
        );

    \I__5000\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20708\
        );

    \I__4999\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20708\
        );

    \I__4998\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20705\
        );

    \I__4997\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20702\
        );

    \I__4996\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20699\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__20734\,
            I => \N__20694\
        );

    \I__4994\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20689\
        );

    \I__4993\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20689\
        );

    \I__4992\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20686\
        );

    \I__4991\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20683\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20680\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20677\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20672\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20672\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__20713\,
            I => \N__20667\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__20708\,
            I => \N__20662\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20662\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__20702\,
            I => \N__20657\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20657\
        );

    \I__4981\ : InMux
    port map (
            O => \N__20698\,
            I => \N__20654\
        );

    \I__4980\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20651\
        );

    \I__4979\ : Span4Mux_s2_h
    port map (
            O => \N__20694\,
            I => \N__20648\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__20689\,
            I => \N__20641\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__20686\,
            I => \N__20641\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20641\
        );

    \I__4975\ : Span4Mux_v
    port map (
            O => \N__20680\,
            I => \N__20634\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__20677\,
            I => \N__20634\
        );

    \I__4973\ : Span4Mux_s3_h
    port map (
            O => \N__20672\,
            I => \N__20634\
        );

    \I__4972\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20629\
        );

    \I__4971\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20629\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__20667\,
            I => bu_rx_data_2
        );

    \I__4969\ : Odrv12
    port map (
            O => \N__20662\,
            I => bu_rx_data_2
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__20657\,
            I => bu_rx_data_2
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__20654\,
            I => bu_rx_data_2
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__20651\,
            I => bu_rx_data_2
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__20648\,
            I => bu_rx_data_2
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__20641\,
            I => bu_rx_data_2
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__20634\,
            I => bu_rx_data_2
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__20629\,
            I => bu_rx_data_2
        );

    \I__4961\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20605\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \N__20599\
        );

    \I__4959\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20596\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20591\
        );

    \I__4957\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20588\
        );

    \I__4956\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20585\
        );

    \I__4955\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20582\
        );

    \I__4954\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20579\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__20596\,
            I => \N__20574\
        );

    \I__4952\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20565\
        );

    \I__4951\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20565\
        );

    \I__4950\ : Span4Mux_v
    port map (
            O => \N__20591\,
            I => \N__20558\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20558\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20558\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20553\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__20579\,
            I => \N__20553\
        );

    \I__4945\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20548\
        );

    \I__4944\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20548\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__20574\,
            I => \N__20545\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20542\
        );

    \I__4941\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20537\
        );

    \I__4940\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20537\
        );

    \I__4939\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20534\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__20565\,
            I => \N__20531\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__20558\,
            I => \N__20528\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__20553\,
            I => \N__20525\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__20548\,
            I => bu_rx_data_5
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__20545\,
            I => bu_rx_data_5
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__20542\,
            I => bu_rx_data_5
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20537\,
            I => bu_rx_data_5
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__20534\,
            I => bu_rx_data_5
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__20531\,
            I => bu_rx_data_5
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__20528\,
            I => bu_rx_data_5
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__20525\,
            I => bu_rx_data_5
        );

    \I__4927\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20503\
        );

    \I__4926\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20500\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__20506\,
            I => \N__20493\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__20503\,
            I => \N__20483\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20483\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20478\
        );

    \I__4921\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20478\
        );

    \I__4920\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20473\
        );

    \I__4919\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20473\
        );

    \I__4918\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20468\
        );

    \I__4917\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20465\
        );

    \I__4916\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20462\
        );

    \I__4915\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20459\
        );

    \I__4914\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20454\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20454\
        );

    \I__4912\ : Span4Mux_s2_v
    port map (
            O => \N__20483\,
            I => \N__20451\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__20478\,
            I => \N__20448\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20445\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20472\,
            I => \N__20440\
        );

    \I__4908\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20440\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20437\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20432\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20432\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__20459\,
            I => \N__20429\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20423\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__20451\,
            I => \N__20418\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__20448\,
            I => \N__20418\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__20445\,
            I => \N__20411\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__20440\,
            I => \N__20411\
        );

    \I__4898\ : Span4Mux_s2_h
    port map (
            O => \N__20437\,
            I => \N__20411\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__20432\,
            I => \N__20406\
        );

    \I__4896\ : Span4Mux_s2_h
    port map (
            O => \N__20429\,
            I => \N__20406\
        );

    \I__4895\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20399\
        );

    \I__4894\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20399\
        );

    \I__4893\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20399\
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__20423\,
            I => bu_rx_data_3
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__20418\,
            I => bu_rx_data_3
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__20411\,
            I => bu_rx_data_3
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__20406\,
            I => bu_rx_data_3
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__20399\,
            I => bu_rx_data_3
        );

    \I__4887\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20381\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20381\
        );

    \I__4885\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20376\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__20381\,
            I => \N__20370\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20367\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20364\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20376\,
            I => \N__20359\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20356\
        );

    \I__4879\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20353\
        );

    \I__4878\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20350\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__20370\,
            I => \N__20347\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20344\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__20364\,
            I => \N__20341\
        );

    \I__4874\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20336\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20336\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__20359\,
            I => \N__20331\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20331\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__20353\,
            I => \N__20328\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__20350\,
            I => \N__20325\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__20347\,
            I => \N__20320\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__20344\,
            I => \N__20320\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__20341\,
            I => \N__20317\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__20336\,
            I => bu_rx_data_7
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__20331\,
            I => bu_rx_data_7
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__20328\,
            I => bu_rx_data_7
        );

    \I__4862\ : Odrv12
    port map (
            O => \N__20325\,
            I => bu_rx_data_7
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__20320\,
            I => bu_rx_data_7
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__20317\,
            I => bu_rx_data_7
        );

    \I__4859\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20299\
        );

    \I__4858\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20292\
        );

    \I__4857\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20289\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20281\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20278\
        );

    \I__4854\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20273\
        );

    \I__4853\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20273\
        );

    \I__4852\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20270\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20265\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20265\
        );

    \I__4849\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20258\
        );

    \I__4848\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20258\
        );

    \I__4847\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20255\
        );

    \I__4846\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20251\
        );

    \I__4845\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20247\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__20281\,
            I => \N__20241\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20241\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__20273\,
            I => \N__20234\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20234\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__20265\,
            I => \N__20234\
        );

    \I__4839\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20229\
        );

    \I__4838\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20229\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20224\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__20255\,
            I => \N__20224\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__20254\,
            I => \N__20220\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20217\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20214\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20211\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20208\
        );

    \I__4830\ : Sp12to4
    port map (
            O => \N__20241\,
            I => \N__20205\
        );

    \I__4829\ : Span4Mux_v
    port map (
            O => \N__20234\,
            I => \N__20200\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__20229\,
            I => \N__20200\
        );

    \I__4827\ : Span4Mux_v
    port map (
            O => \N__20224\,
            I => \N__20197\
        );

    \I__4826\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20194\
        );

    \I__4825\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20191\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__20217\,
            I => \N__20184\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20184\
        );

    \I__4822\ : Span4Mux_s2_h
    port map (
            O => \N__20211\,
            I => \N__20184\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__20208\,
            I => bu_rx_data_1
        );

    \I__4820\ : Odrv12
    port map (
            O => \N__20205\,
            I => bu_rx_data_1
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__20200\,
            I => bu_rx_data_1
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__20197\,
            I => bu_rx_data_1
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__20194\,
            I => bu_rx_data_1
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__20191\,
            I => bu_rx_data_1
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__20184\,
            I => bu_rx_data_1
        );

    \I__4814\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20164\
        );

    \I__4813\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20152\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20149\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20146\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__20163\,
            I => \N__20143\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20139\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20136\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20133\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20130\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20125\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20125\
        );

    \I__4803\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20122\
        );

    \I__4802\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20119\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20152\,
            I => \N__20116\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__20149\,
            I => \N__20113\
        );

    \I__4799\ : Span4Mux_s1_h
    port map (
            O => \N__20146\,
            I => \N__20110\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20107\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20104\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20101\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__20136\,
            I => \N__20098\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20091\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__20130\,
            I => \N__20091\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20091\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20084\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20119\,
            I => \N__20084\
        );

    \I__4789\ : Span4Mux_s3_h
    port map (
            O => \N__20116\,
            I => \N__20084\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__20113\,
            I => \N__20079\
        );

    \I__4787\ : Span4Mux_h
    port map (
            O => \N__20110\,
            I => \N__20079\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__20107\,
            I => \N__20074\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20074\
        );

    \I__4784\ : Span4Mux_s3_h
    port map (
            O => \N__20101\,
            I => \N__20065\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__20098\,
            I => \N__20065\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__20091\,
            I => \N__20065\
        );

    \I__4781\ : Span4Mux_v
    port map (
            O => \N__20084\,
            I => \N__20065\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__20079\,
            I => bu_rx_data_6
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__20074\,
            I => bu_rx_data_6
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__20065\,
            I => bu_rx_data_6
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__20058\,
            I => \N__20053\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20049\
        );

    \I__4775\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20045\
        );

    \I__4774\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20042\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__20052\,
            I => \N__20039\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20034\
        );

    \I__4771\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20031\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20045\,
            I => \N__20026\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__20042\,
            I => \N__20023\
        );

    \I__4768\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20020\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20017\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20014\
        );

    \I__4765\ : Span4Mux_v
    port map (
            O => \N__20034\,
            I => \N__20007\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20007\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20004\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20000\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__20026\,
            I => \N__19993\
        );

    \I__4760\ : Span4Mux_s1_h
    port map (
            O => \N__20023\,
            I => \N__19993\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20020\,
            I => \N__19993\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20017\,
            I => \N__19988\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__19988\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20013\,
            I => \N__19983\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20012\,
            I => \N__19983\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__20007\,
            I => \N__19978\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__19978\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19975\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19970\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__19993\,
            I => \N__19970\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__19988\,
            I => \N__19967\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__19983\,
            I => bu_rx_data_4
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__19978\,
            I => bu_rx_data_4
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__19975\,
            I => bu_rx_data_4
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__19970\,
            I => bu_rx_data_4
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__19967\,
            I => bu_rx_data_4
        );

    \I__4743\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19952\
        );

    \I__4742\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19945\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19942\
        );

    \I__4740\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19937\
        );

    \I__4739\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19937\
        );

    \I__4738\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19934\
        );

    \I__4737\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19930\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19919\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__19942\,
            I => \N__19919\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__19937\,
            I => \N__19919\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19916\
        );

    \I__4732\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19913\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__19930\,
            I => \N__19909\
        );

    \I__4730\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19906\
        );

    \I__4729\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19902\
        );

    \I__4728\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19897\
        );

    \I__4727\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19897\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__19919\,
            I => \N__19892\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__19916\,
            I => \N__19892\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19889\
        );

    \I__4723\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19885\
        );

    \I__4722\ : Span4Mux_s2_v
    port map (
            O => \N__19909\,
            I => \N__19880\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__19906\,
            I => \N__19880\
        );

    \I__4720\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19877\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__19902\,
            I => \N__19874\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19869\
        );

    \I__4717\ : Span4Mux_v
    port map (
            O => \N__19892\,
            I => \N__19864\
        );

    \I__4716\ : Span4Mux_v
    port map (
            O => \N__19889\,
            I => \N__19864\
        );

    \I__4715\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19861\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19858\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__19880\,
            I => \N__19853\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19853\
        );

    \I__4711\ : Span12Mux_s8_v
    port map (
            O => \N__19874\,
            I => \N__19850\
        );

    \I__4710\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19847\
        );

    \I__4709\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19844\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__19869\,
            I => \N__19839\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__19864\,
            I => \N__19839\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__19861\,
            I => \N__19832\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__19858\,
            I => \N__19832\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__19853\,
            I => \N__19832\
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__19850\,
            I => bu_rx_data_0
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__19847\,
            I => bu_rx_data_0
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__19844\,
            I => bu_rx_data_0
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__19839\,
            I => bu_rx_data_0
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__19832\,
            I => bu_rx_data_0
        );

    \I__4698\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__19815\,
            I => \Lab_UT.dictrl.g0_5_o4_3\
        );

    \I__4695\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19806\
        );

    \I__4694\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19803\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__19810\,
            I => \N__19799\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__19809\,
            I => \N__19796\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19788\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19788\
        );

    \I__4689\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19785\
        );

    \I__4688\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19782\
        );

    \I__4687\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19775\
        );

    \I__4686\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19771\
        );

    \I__4685\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19766\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19766\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__19788\,
            I => \N__19763\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19758\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N__19758\
        );

    \I__4680\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19750\
        );

    \I__4679\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19750\
        );

    \I__4678\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19745\
        );

    \I__4677\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19745\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__19775\,
            I => \N__19740\
        );

    \I__4675\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19736\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19727\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19727\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__19763\,
            I => \N__19727\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__19758\,
            I => \N__19727\
        );

    \I__4670\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19724\
        );

    \I__4669\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19721\
        );

    \I__4668\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19718\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19713\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19713\
        );

    \I__4665\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19708\
        );

    \I__4664\ : InMux
    port map (
            O => \N__19743\,
            I => \N__19708\
        );

    \I__4663\ : Span4Mux_v
    port map (
            O => \N__19740\,
            I => \N__19705\
        );

    \I__4662\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19702\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19695\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19695\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19695\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__19721\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__19718\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__19713\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__19708\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__19705\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__19702\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__19695\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__19680\,
            I => \Lab_UT.dictrl.g0_5_o4_4_cascade_\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__19677\,
            I => \N__19673\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19666\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19662\
        );

    \I__4647\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19659\
        );

    \I__4646\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19656\
        );

    \I__4645\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19651\
        );

    \I__4644\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19642\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19666\,
            I => \N__19638\
        );

    \I__4642\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19635\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19632\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__19659\,
            I => \N__19629\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__19656\,
            I => \N__19626\
        );

    \I__4638\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19621\
        );

    \I__4637\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19621\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__19651\,
            I => \N__19618\
        );

    \I__4635\ : InMux
    port map (
            O => \N__19650\,
            I => \N__19615\
        );

    \I__4634\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19612\
        );

    \I__4633\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19609\
        );

    \I__4632\ : InMux
    port map (
            O => \N__19647\,
            I => \N__19604\
        );

    \I__4631\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19604\
        );

    \I__4630\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19601\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__19642\,
            I => \N__19598\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19595\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__19638\,
            I => \N__19590\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19590\
        );

    \I__4625\ : Span4Mux_s3_h
    port map (
            O => \N__19632\,
            I => \N__19585\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__19629\,
            I => \N__19585\
        );

    \I__4623\ : Span4Mux_v
    port map (
            O => \N__19626\,
            I => \N__19578\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19578\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__19618\,
            I => \N__19578\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__19615\,
            I => \N__19569\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__19612\,
            I => \N__19569\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__19609\,
            I => \N__19569\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19604\,
            I => \N__19569\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19601\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__19598\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__19595\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__19590\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__19585\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__19578\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__19569\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__19548\,
            I => \Lab_UT.dictrl.N_11\
        );

    \I__4606\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19542\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__19539\,
            I => \buart.Z_rx.P7_mux\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N_16_mux\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__19530\,
            I => \shifter_7_rep1_RNIG7Q01_cascade_\
        );

    \I__4600\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__19521\,
            I => \N__19517\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19514\
        );

    \I__4596\ : Span4Mux_s3_h
    port map (
            O => \N__19517\,
            I => \N__19509\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19509\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__19506\,
            I => \N_97\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__19500\,
            I => \N__19492\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19489\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19486\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19483\
        );

    \I__4587\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19480\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19477\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__19492\,
            I => \N__19472\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19472\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19486\,
            I => \N__19469\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19466\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19461\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19461\
        );

    \I__4579\ : Span4Mux_h
    port map (
            O => \N__19472\,
            I => \N__19458\
        );

    \I__4578\ : Sp12to4
    port map (
            O => \N__19469\,
            I => \N__19455\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__19466\,
            I => \N__19452\
        );

    \I__4576\ : Span4Mux_h
    port map (
            O => \N__19461\,
            I => \N__19449\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__19458\,
            I => \N__19446\
        );

    \I__4574\ : Odrv12
    port map (
            O => \N__19455\,
            I => bu_rx_data_4_rep1
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__19452\,
            I => bu_rx_data_4_rep1
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__19449\,
            I => bu_rx_data_4_rep1
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__19446\,
            I => bu_rx_data_4_rep1
        );

    \I__4570\ : IoInMux
    port map (
            O => \N__19437\,
            I => \N__19434\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__19431\,
            I => bu_rx_data_rdy_0
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__19428\,
            I => \N__19425\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19414\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19409\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19409\
        );

    \I__4562\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19404\
        );

    \I__4561\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19397\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19397\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__19414\,
            I => \N__19390\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19390\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19385\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19385\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19382\
        );

    \I__4554\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19377\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19377\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__19397\,
            I => \N__19373\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19370\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19367\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__19390\,
            I => \N__19362\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N__19362\
        );

    \I__4547\ : Span4Mux_v
    port map (
            O => \N__19382\,
            I => \N__19357\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__19377\,
            I => \N__19357\
        );

    \I__4545\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19354\
        );

    \I__4544\ : Span12Mux_s6_v
    port map (
            O => \N__19373\,
            I => \N__19351\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19370\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19367\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__19362\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__19357\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19354\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4538\ : Odrv12
    port map (
            O => \N__19351\,
            I => \Lab_UT_dictrl_state_3_rep2\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__19338\,
            I => \Lab_UT.dictrl.g0_5_a4_1_5_cascade_\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \Lab_UT.dictrl.N_13_cascade_\
        );

    \I__4535\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__19326\,
            I => \N__19323\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__19323\,
            I => \Lab_UT.dictrl.N_90\
        );

    \I__4531\ : CEMux
    port map (
            O => \N__19320\,
            I => \N__19296\
        );

    \I__4530\ : CEMux
    port map (
            O => \N__19319\,
            I => \N__19296\
        );

    \I__4529\ : CEMux
    port map (
            O => \N__19318\,
            I => \N__19296\
        );

    \I__4528\ : CEMux
    port map (
            O => \N__19317\,
            I => \N__19296\
        );

    \I__4527\ : CEMux
    port map (
            O => \N__19316\,
            I => \N__19296\
        );

    \I__4526\ : CEMux
    port map (
            O => \N__19315\,
            I => \N__19296\
        );

    \I__4525\ : CEMux
    port map (
            O => \N__19314\,
            I => \N__19296\
        );

    \I__4524\ : CEMux
    port map (
            O => \N__19313\,
            I => \N__19296\
        );

    \I__4523\ : GlobalMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__4522\ : gio2CtrlBuf
    port map (
            O => \N__19293\,
            I => \buart.Z_rx.sample_g\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__19290\,
            I => \N__19279\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19275\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19272\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19269\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19266\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19263\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19260\
        );

    \I__4514\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19257\
        );

    \I__4513\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19254\
        );

    \I__4512\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19251\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19248\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19245\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19242\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19196\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__19266\,
            I => \N__19193\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__19263\,
            I => \N__19190\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__19260\,
            I => \N__19187\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19184\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19181\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19251\,
            I => \N__19163\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19160\
        );

    \I__4500\ : Glb2LocalMux
    port map (
            O => \N__19245\,
            I => \N__19023\
        );

    \I__4499\ : Glb2LocalMux
    port map (
            O => \N__19242\,
            I => \N__19023\
        );

    \I__4498\ : SRMux
    port map (
            O => \N__19241\,
            I => \N__19023\
        );

    \I__4497\ : SRMux
    port map (
            O => \N__19240\,
            I => \N__19023\
        );

    \I__4496\ : SRMux
    port map (
            O => \N__19239\,
            I => \N__19023\
        );

    \I__4495\ : SRMux
    port map (
            O => \N__19238\,
            I => \N__19023\
        );

    \I__4494\ : SRMux
    port map (
            O => \N__19237\,
            I => \N__19023\
        );

    \I__4493\ : SRMux
    port map (
            O => \N__19236\,
            I => \N__19023\
        );

    \I__4492\ : SRMux
    port map (
            O => \N__19235\,
            I => \N__19023\
        );

    \I__4491\ : SRMux
    port map (
            O => \N__19234\,
            I => \N__19023\
        );

    \I__4490\ : SRMux
    port map (
            O => \N__19233\,
            I => \N__19023\
        );

    \I__4489\ : SRMux
    port map (
            O => \N__19232\,
            I => \N__19023\
        );

    \I__4488\ : SRMux
    port map (
            O => \N__19231\,
            I => \N__19023\
        );

    \I__4487\ : SRMux
    port map (
            O => \N__19230\,
            I => \N__19023\
        );

    \I__4486\ : SRMux
    port map (
            O => \N__19229\,
            I => \N__19023\
        );

    \I__4485\ : SRMux
    port map (
            O => \N__19228\,
            I => \N__19023\
        );

    \I__4484\ : SRMux
    port map (
            O => \N__19227\,
            I => \N__19023\
        );

    \I__4483\ : SRMux
    port map (
            O => \N__19226\,
            I => \N__19023\
        );

    \I__4482\ : SRMux
    port map (
            O => \N__19225\,
            I => \N__19023\
        );

    \I__4481\ : SRMux
    port map (
            O => \N__19224\,
            I => \N__19023\
        );

    \I__4480\ : SRMux
    port map (
            O => \N__19223\,
            I => \N__19023\
        );

    \I__4479\ : SRMux
    port map (
            O => \N__19222\,
            I => \N__19023\
        );

    \I__4478\ : SRMux
    port map (
            O => \N__19221\,
            I => \N__19023\
        );

    \I__4477\ : SRMux
    port map (
            O => \N__19220\,
            I => \N__19023\
        );

    \I__4476\ : SRMux
    port map (
            O => \N__19219\,
            I => \N__19023\
        );

    \I__4475\ : SRMux
    port map (
            O => \N__19218\,
            I => \N__19023\
        );

    \I__4474\ : SRMux
    port map (
            O => \N__19217\,
            I => \N__19023\
        );

    \I__4473\ : SRMux
    port map (
            O => \N__19216\,
            I => \N__19023\
        );

    \I__4472\ : SRMux
    port map (
            O => \N__19215\,
            I => \N__19023\
        );

    \I__4471\ : SRMux
    port map (
            O => \N__19214\,
            I => \N__19023\
        );

    \I__4470\ : SRMux
    port map (
            O => \N__19213\,
            I => \N__19023\
        );

    \I__4469\ : SRMux
    port map (
            O => \N__19212\,
            I => \N__19023\
        );

    \I__4468\ : SRMux
    port map (
            O => \N__19211\,
            I => \N__19023\
        );

    \I__4467\ : SRMux
    port map (
            O => \N__19210\,
            I => \N__19023\
        );

    \I__4466\ : SRMux
    port map (
            O => \N__19209\,
            I => \N__19023\
        );

    \I__4465\ : SRMux
    port map (
            O => \N__19208\,
            I => \N__19023\
        );

    \I__4464\ : SRMux
    port map (
            O => \N__19207\,
            I => \N__19023\
        );

    \I__4463\ : SRMux
    port map (
            O => \N__19206\,
            I => \N__19023\
        );

    \I__4462\ : SRMux
    port map (
            O => \N__19205\,
            I => \N__19023\
        );

    \I__4461\ : SRMux
    port map (
            O => \N__19204\,
            I => \N__19023\
        );

    \I__4460\ : SRMux
    port map (
            O => \N__19203\,
            I => \N__19023\
        );

    \I__4459\ : SRMux
    port map (
            O => \N__19202\,
            I => \N__19023\
        );

    \I__4458\ : SRMux
    port map (
            O => \N__19201\,
            I => \N__19023\
        );

    \I__4457\ : SRMux
    port map (
            O => \N__19200\,
            I => \N__19023\
        );

    \I__4456\ : SRMux
    port map (
            O => \N__19199\,
            I => \N__19023\
        );

    \I__4455\ : Glb2LocalMux
    port map (
            O => \N__19196\,
            I => \N__19023\
        );

    \I__4454\ : Glb2LocalMux
    port map (
            O => \N__19193\,
            I => \N__19023\
        );

    \I__4453\ : Glb2LocalMux
    port map (
            O => \N__19190\,
            I => \N__19023\
        );

    \I__4452\ : Glb2LocalMux
    port map (
            O => \N__19187\,
            I => \N__19023\
        );

    \I__4451\ : Glb2LocalMux
    port map (
            O => \N__19184\,
            I => \N__19023\
        );

    \I__4450\ : Glb2LocalMux
    port map (
            O => \N__19181\,
            I => \N__19023\
        );

    \I__4449\ : SRMux
    port map (
            O => \N__19180\,
            I => \N__19023\
        );

    \I__4448\ : SRMux
    port map (
            O => \N__19179\,
            I => \N__19023\
        );

    \I__4447\ : SRMux
    port map (
            O => \N__19178\,
            I => \N__19023\
        );

    \I__4446\ : SRMux
    port map (
            O => \N__19177\,
            I => \N__19023\
        );

    \I__4445\ : SRMux
    port map (
            O => \N__19176\,
            I => \N__19023\
        );

    \I__4444\ : SRMux
    port map (
            O => \N__19175\,
            I => \N__19023\
        );

    \I__4443\ : SRMux
    port map (
            O => \N__19174\,
            I => \N__19023\
        );

    \I__4442\ : SRMux
    port map (
            O => \N__19173\,
            I => \N__19023\
        );

    \I__4441\ : SRMux
    port map (
            O => \N__19172\,
            I => \N__19023\
        );

    \I__4440\ : SRMux
    port map (
            O => \N__19171\,
            I => \N__19023\
        );

    \I__4439\ : SRMux
    port map (
            O => \N__19170\,
            I => \N__19023\
        );

    \I__4438\ : SRMux
    port map (
            O => \N__19169\,
            I => \N__19023\
        );

    \I__4437\ : SRMux
    port map (
            O => \N__19168\,
            I => \N__19023\
        );

    \I__4436\ : SRMux
    port map (
            O => \N__19167\,
            I => \N__19023\
        );

    \I__4435\ : SRMux
    port map (
            O => \N__19166\,
            I => \N__19023\
        );

    \I__4434\ : Glb2LocalMux
    port map (
            O => \N__19163\,
            I => \N__19023\
        );

    \I__4433\ : Glb2LocalMux
    port map (
            O => \N__19160\,
            I => \N__19023\
        );

    \I__4432\ : GlobalMux
    port map (
            O => \N__19023\,
            I => \N__19020\
        );

    \I__4431\ : gio2CtrlBuf
    port map (
            O => \N__19020\,
            I => rst_g
        );

    \I__4430\ : InMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__4428\ : Span4Mux_v
    port map (
            O => \N__19011\,
            I => \N__19006\
        );

    \I__4427\ : InMux
    port map (
            O => \N__19010\,
            I => \N__19003\
        );

    \I__4426\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19000\
        );

    \I__4425\ : IoSpan4Mux
    port map (
            O => \N__19006\,
            I => \N__18994\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19003\,
            I => \N__18994\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19000\,
            I => \N__18991\
        );

    \I__4422\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18988\
        );

    \I__4421\ : Span4Mux_s2_h
    port map (
            O => \N__18994\,
            I => \N__18983\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__18991\,
            I => \N__18980\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__18988\,
            I => \N__18977\
        );

    \I__4418\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18972\
        );

    \I__4417\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18972\
        );

    \I__4416\ : Span4Mux_h
    port map (
            O => \N__18983\,
            I => \N__18969\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__18980\,
            I => bu_rx_data_rdy
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__18977\,
            I => bu_rx_data_rdy
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__18972\,
            I => bu_rx_data_rdy
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__18969\,
            I => bu_rx_data_rdy
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__18960\,
            I => \N__18957\
        );

    \I__4410\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18954\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__4408\ : Span4Mux_s1_h
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__18948\,
            I => \Lab_UT.dictrl.m25Z0Z_0\
        );

    \I__4406\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18937\
        );

    \I__4405\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18932\
        );

    \I__4404\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18932\
        );

    \I__4403\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18927\
        );

    \I__4402\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18927\
        );

    \I__4401\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18924\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18917\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18917\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__18927\,
            I => \N__18917\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__18924\,
            I => bu_rx_data_fast_2
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__18917\,
            I => bu_rx_data_fast_2
        );

    \I__4395\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18905\
        );

    \I__4394\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18905\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__18910\,
            I => \N__18902\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18896\
        );

    \I__4391\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18893\
        );

    \I__4390\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18886\
        );

    \I__4389\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18886\
        );

    \I__4388\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18886\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__18896\,
            I => \N__18879\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18879\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__18886\,
            I => \N__18879\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__18879\,
            I => \buart__rx_shifter_fast_5\
        );

    \I__4383\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18869\
        );

    \I__4382\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18869\
        );

    \I__4381\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18863\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18860\
        );

    \I__4379\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18855\
        );

    \I__4378\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18855\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__18866\,
            I => \N__18847\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__18863\,
            I => \N__18843\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__18860\,
            I => \N__18838\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__18855\,
            I => \N__18838\
        );

    \I__4373\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18833\
        );

    \I__4372\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18833\
        );

    \I__4371\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18830\
        );

    \I__4370\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18827\
        );

    \I__4369\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18820\
        );

    \I__4368\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18820\
        );

    \I__4367\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18820\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__18843\,
            I => \N__18817\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__18838\,
            I => \N__18814\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18811\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__18830\,
            I => bu_rx_data_2_rep1
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__18827\,
            I => bu_rx_data_2_rep1
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__18820\,
            I => bu_rx_data_2_rep1
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__18817\,
            I => bu_rx_data_2_rep1
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__18814\,
            I => bu_rx_data_2_rep1
        );

    \I__4358\ : Odrv12
    port map (
            O => \N__18811\,
            I => bu_rx_data_2_rep1
        );

    \I__4357\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18795\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__4355\ : Span4Mux_s3_h
    port map (
            O => \N__18792\,
            I => \N__18783\
        );

    \I__4354\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18780\
        );

    \I__4353\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18777\
        );

    \I__4352\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18772\
        );

    \I__4351\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18772\
        );

    \I__4350\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18767\
        );

    \I__4349\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18767\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__18783\,
            I => \Lab_UT.dictrl.N_103_mux\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__18780\,
            I => \Lab_UT.dictrl.N_103_mux\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__18777\,
            I => \Lab_UT.dictrl.N_103_mux\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18772\,
            I => \Lab_UT.dictrl.N_103_mux\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__18767\,
            I => \Lab_UT.dictrl.N_103_mux\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__18756\,
            I => \Lab_UT.dictrl.N_4_0_cascade_\
        );

    \I__4342\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18744\
        );

    \I__4341\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18739\
        );

    \I__4340\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18739\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__18750\,
            I => \N__18735\
        );

    \I__4338\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18730\
        );

    \I__4337\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18730\
        );

    \I__4336\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18727\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__18744\,
            I => \N__18724\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__18739\,
            I => \N__18721\
        );

    \I__4333\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18716\
        );

    \I__4332\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18713\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18710\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18703\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__18724\,
            I => \N__18703\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__18721\,
            I => \N__18703\
        );

    \I__4327\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18698\
        );

    \I__4326\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18698\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__18716\,
            I => \N__18695\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__18713\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__18710\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__18703\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__18698\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__4320\ : Odrv12
    port map (
            O => \N__18695\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__4319\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18681\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__18675\,
            I => \Lab_UT.dictrl.N_12_0\
        );

    \I__4315\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__18669\,
            I => \N__18666\
        );

    \I__4313\ : Odrv12
    port map (
            O => \N__18666\,
            I => \Lab_UT.LdASones\
        );

    \I__4312\ : CEMux
    port map (
            O => \N__18663\,
            I => \N__18659\
        );

    \I__4311\ : CEMux
    port map (
            O => \N__18662\,
            I => \N__18656\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__18659\,
            I => \N__18653\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__18656\,
            I => \N__18650\
        );

    \I__4308\ : Sp12to4
    port map (
            O => \N__18653\,
            I => \N__18647\
        );

    \I__4307\ : Span4Mux_v
    port map (
            O => \N__18650\,
            I => \N__18644\
        );

    \I__4306\ : Span12Mux_v
    port map (
            O => \N__18647\,
            I => \N__18641\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__4304\ : Odrv12
    port map (
            O => \N__18641\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__18638\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__18633\,
            I => \N__18629\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__18632\,
            I => \N__18624\
        );

    \I__4300\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18621\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__18628\,
            I => \N__18618\
        );

    \I__4298\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18615\
        );

    \I__4297\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18612\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__18621\,
            I => \N__18609\
        );

    \I__4295\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18606\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__18615\,
            I => \N__18602\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__18612\,
            I => \N__18599\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__18609\,
            I => \N__18594\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18594\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__18605\,
            I => \N__18591\
        );

    \I__4289\ : Span12Mux_s5_h
    port map (
            O => \N__18602\,
            I => \N__18588\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__18599\,
            I => \N__18585\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__18594\,
            I => \N__18582\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18579\
        );

    \I__4285\ : Odrv12
    port map (
            O => \N__18588\,
            I => bu_rx_data_7_rep1
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__18585\,
            I => bu_rx_data_7_rep1
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__18582\,
            I => bu_rx_data_7_rep1
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18579\,
            I => bu_rx_data_7_rep1
        );

    \I__4281\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__18567\,
            I => \shifter_7_rep1_RNIG7Q01\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__18564\,
            I => \Lab_UT.dictrl.N_77_cascade_\
        );

    \I__4278\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__18555\,
            I => \Lab_UT.dictrl.m73Z0Z_1\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18549\,
            I => \Lab_UT.dictrl.m77_ns_1\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__18546\,
            I => \Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_\
        );

    \I__4272\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18539\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18536\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18533\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18530\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__18533\,
            I => \N__18527\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__18530\,
            I => \Lab_UT.dictrl.i9_mux_0_0\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__18527\,
            I => \Lab_UT.dictrl.i9_mux_0_0\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18516\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18516\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18512\
        );

    \I__4262\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18509\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__18512\,
            I => \Lab_UT.dictrl.N_106_mux\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__18509\,
            I => \Lab_UT.dictrl.N_106_mux\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18498\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__18498\,
            I => \Lab_UT.dictrl.m51_0\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18495\,
            I => \N__18490\
        );

    \I__4255\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18487\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18484\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18490\,
            I => \N__18481\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18478\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__18484\,
            I => \N__18472\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__18481\,
            I => \N__18472\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__18478\,
            I => \N__18469\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__18477\,
            I => \N__18466\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__18472\,
            I => \N__18461\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__18469\,
            I => \N__18461\
        );

    \I__4245\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18458\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__18461\,
            I => \Lab_UT.dictrl.state_i_3_1\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18458\,
            I => \Lab_UT.dictrl.state_i_3_1\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__18453\,
            I => \Lab_UT.dictrl.N_118_mux_cascade_\
        );

    \I__4241\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18447\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18447\,
            I => \N__18444\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__18444\,
            I => \Lab_UT.dictrl.next_state_latmux_3_1_1\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18438\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18438\,
            I => \N__18435\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__18435\,
            I => \N__18432\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__18432\,
            I => \Lab_UT.dictrl.g0_17_a6_3Z0Z_7\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__18429\,
            I => \N__18425\
        );

    \I__4233\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18420\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18414\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18414\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18411\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18408\
        );

    \I__4228\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18405\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__18414\,
            I => \N__18402\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__18411\,
            I => \N__18399\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__18408\,
            I => \N__18396\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__18405\,
            I => \N__18391\
        );

    \I__4223\ : Span4Mux_h
    port map (
            O => \N__18402\,
            I => \N__18391\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__18399\,
            I => \buart__rx_shifter_fast_0\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18396\,
            I => \buart__rx_shifter_fast_0\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__18391\,
            I => \buart__rx_shifter_fast_0\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__18384\,
            I => \N__18376\
        );

    \I__4218\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18370\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18370\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18365\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18365\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18362\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18359\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18356\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18348\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18348\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18362\,
            I => \N__18343\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__18359\,
            I => \N__18343\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__18356\,
            I => \N__18340\
        );

    \I__4206\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18337\
        );

    \I__4205\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18332\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18332\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__18348\,
            I => \N__18329\
        );

    \I__4202\ : Span4Mux_s3_h
    port map (
            O => \N__18343\,
            I => \N__18326\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__18340\,
            I => bu_rx_data_1_rep1
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18337\,
            I => bu_rx_data_1_rep1
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__18332\,
            I => bu_rx_data_1_rep1
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__18329\,
            I => bu_rx_data_1_rep1
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__18326\,
            I => bu_rx_data_1_rep1
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__18315\,
            I => \N__18311\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18303\
        );

    \I__4194\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18303\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18303\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__18303\,
            I => \N__18299\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18294\
        );

    \I__4190\ : Span4Mux_v
    port map (
            O => \N__18299\,
            I => \N__18291\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__18298\,
            I => \N__18288\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18283\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18294\,
            I => \N__18278\
        );

    \I__4186\ : Sp12to4
    port map (
            O => \N__18291\,
            I => \N__18278\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18271\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18271\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18271\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__18283\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4181\ : Odrv12
    port map (
            O => \N__18278\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__18271\,
            I => \Lab_UT.dictrl.next_state_1_3\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18261\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__18261\,
            I => \Lab_UT.dictrl.P6_mux_0\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__18258\,
            I => \N__18254\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18250\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18247\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18244\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18250\,
            I => \N__18241\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__18247\,
            I => \N__18238\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__18244\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__18241\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__18238\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__18231\,
            I => \N__18228\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18222\,
            I => \Lab_UT.dictrl.N_114_mux\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18216\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18216\,
            I => \Lab_UT.dictrl.N_69\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__18213\,
            I => \N__18209\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18204\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18204\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18204\,
            I => \Lab_UT.dictrl.i10_mux\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__18201\,
            I => \Lab_UT.dictrl.N_69_cascade_\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18192\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__18192\,
            I => \N__18189\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__18189\,
            I => \Lab_UT.dictrl.next_state_1_0_3\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18183\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18180\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__18180\,
            I => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__18177\,
            I => \N__18171\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \N__18168\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18165\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18158\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18158\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18158\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18155\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__18158\,
            I => \N__18150\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18155\,
            I => \N__18150\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__18150\,
            I => \N__18147\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__18147\,
            I => \Lab_UT.dictrl.g0_17_a6_0_1\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18138\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18138\,
            I => \Lab_UT.dictrl.P6_mux\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18128\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18128\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18125\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18128\,
            I => \N__18122\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18125\,
            I => \N__18119\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__18122\,
            I => \N__18116\
        );

    \I__4130\ : Span4Mux_h
    port map (
            O => \N__18119\,
            I => \N__18113\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__18116\,
            I => \Lab_UT.dictrl.N_189\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__18113\,
            I => \Lab_UT.dictrl.N_189\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18098\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18098\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18095\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18098\,
            I => \Lab_UT.dictrl.m40_N_5_mux\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18095\,
            I => \Lab_UT.dictrl.m40_N_5_mux\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18086\
        );

    \I__4120\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18083\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18086\,
            I => \Lab_UT.dictrl.N_77\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__18083\,
            I => \Lab_UT.dictrl.N_77\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18072\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18072\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18072\,
            I => \Lab_UT.dictrl.alarmstate8Z0Z_4\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18065\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \N__18062\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18057\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18054\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18051\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18048\
        );

    \I__4108\ : Span4Mux_s3_h
    port map (
            O => \N__18057\,
            I => \N__18041\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18041\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18051\,
            I => \N__18036\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18048\,
            I => \N__18036\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18029\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18029\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__18041\,
            I => \N__18026\
        );

    \I__4101\ : Span4Mux_v
    port map (
            O => \N__18036\,
            I => \N__18023\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18020\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18017\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18029\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__18026\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__18023\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18020\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18017\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18006\,
            I => \N__18003\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17999\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__18002\,
            I => \N__17995\
        );

    \I__4090\ : Span4Mux_h
    port map (
            O => \N__17999\,
            I => \N__17991\
        );

    \I__4089\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17988\
        );

    \I__4088\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17985\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__17994\,
            I => \N__17982\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__17991\,
            I => \N__17977\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__17988\,
            I => \N__17977\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__17985\,
            I => \N__17974\
        );

    \I__4083\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17971\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__17977\,
            I => \Lab_UT.LdSones\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__17974\,
            I => \Lab_UT.LdSones\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__17971\,
            I => \Lab_UT.LdSones\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17961\,
            I => \N__17957\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__17960\,
            I => \N__17953\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__17957\,
            I => \N__17946\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__17956\,
            I => \N__17943\
        );

    \I__4074\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17940\
        );

    \I__4073\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17937\
        );

    \I__4072\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17932\
        );

    \I__4071\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17932\
        );

    \I__4070\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17929\
        );

    \I__4069\ : Span4Mux_s3_h
    port map (
            O => \N__17946\,
            I => \N__17926\
        );

    \I__4068\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17923\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__17940\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__17937\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__17932\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__17929\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__17926\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__17923\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__4061\ : InMux
    port map (
            O => \N__17910\,
            I => \N__17907\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__17907\,
            I => \Lab_UT.didp.countrce1.q_5_1\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__17904\,
            I => \Lab_UT.dictrl.N_4_cascade_\
        );

    \I__4058\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17898\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__17898\,
            I => \N__17892\
        );

    \I__4056\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17885\
        );

    \I__4055\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17885\
        );

    \I__4054\ : InMux
    port map (
            O => \N__17895\,
            I => \N__17885\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__17892\,
            I => \N__17882\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__17885\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__17882\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__4050\ : InMux
    port map (
            O => \N__17877\,
            I => \N__17873\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__17876\,
            I => \N__17870\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17867\
        );

    \I__4047\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17864\
        );

    \I__4046\ : Odrv12
    port map (
            O => \N__17867\,
            I => \Lab_UT.dictrl.N_81\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__17864\,
            I => \Lab_UT.dictrl.N_81\
        );

    \I__4044\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17856\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__17856\,
            I => \Lab_UT.dictrl.next_state_i_1_2\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__17853\,
            I => \N__17850\
        );

    \I__4041\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17847\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__4038\ : Span4Mux_v
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__4037\ : Odrv4
    port map (
            O => \N__17838\,
            I => \Lab_UT.dictrl.P8_mux\
        );

    \I__4036\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17831\
        );

    \I__4035\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17828\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17821\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17816\
        );

    \I__4032\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17810\
        );

    \I__4031\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17807\
        );

    \I__4030\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17802\
        );

    \I__4029\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17802\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__17821\,
            I => \N__17799\
        );

    \I__4027\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17794\
        );

    \I__4026\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17794\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__17816\,
            I => \N__17791\
        );

    \I__4024\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17784\
        );

    \I__4023\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17784\
        );

    \I__4022\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17784\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__17810\,
            I => \G_183\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__17807\,
            I => \G_183\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__17802\,
            I => \G_183\
        );

    \I__4018\ : Odrv4
    port map (
            O => \N__17799\,
            I => \G_183\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__17794\,
            I => \G_183\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__17791\,
            I => \G_183\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__17784\,
            I => \G_183\
        );

    \I__4014\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17764\
        );

    \I__4013\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17758\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17767\,
            I => \N__17752\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__17764\,
            I => \N__17749\
        );

    \I__4010\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17742\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17742\
        );

    \I__4008\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17742\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17739\
        );

    \I__4006\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17731\
        );

    \I__4005\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17731\
        );

    \I__4004\ : InMux
    port map (
            O => \N__17755\,
            I => \N__17728\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__17752\,
            I => \N__17719\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__17749\,
            I => \N__17719\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17719\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__17739\,
            I => \N__17719\
        );

    \I__3999\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17712\
        );

    \I__3998\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17712\
        );

    \I__3997\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17712\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__17731\,
            I => \G_185\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__17728\,
            I => \G_185\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__17719\,
            I => \G_185\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__17712\,
            I => \G_185\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__17703\,
            I => \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\
        );

    \I__3991\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17697\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__17697\,
            I => \Lab_UT.dictrl.m3_0\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__17694\,
            I => \Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17688\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__17688\,
            I => \G_188\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17682\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__17682\,
            I => \Lab_UT.dictrl.alarmstate8Z0Z_3\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__17679\,
            I => \G_188_cascade_\
        );

    \I__3983\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17673\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__17673\,
            I => \G_187\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__17670\,
            I => \N__17666\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17661\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17661\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__17661\,
            I => \N__17658\
        );

    \I__3977\ : Odrv12
    port map (
            O => \N__17658\,
            I => \G_186\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__17655\,
            I => \G_187_cascade_\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17652\,
            I => \N__17643\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17643\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17643\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__17643\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\
        );

    \I__3971\ : InMux
    port map (
            O => \N__17640\,
            I => \N__17637\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17637\,
            I => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17634\,
            I => \N__17625\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17616\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17616\
        );

    \I__3966\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17616\
        );

    \I__3965\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17616\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__17629\,
            I => \N__17613\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__17628\,
            I => \N__17610\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17607\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17616\,
            I => \N__17604\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17601\
        );

    \I__3959\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17598\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__17607\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__17604\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17601\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17598\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__17589\,
            I => \Lab_UT.dictrl.g0_2Z0Z_2_cascade_\
        );

    \I__3953\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17583\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17583\,
            I => \N__17580\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__17580\,
            I => \Lab_UT.dictrl.m40_N_5_mux_1\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17574\,
            I => \N__17570\
        );

    \I__3948\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17567\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__17570\,
            I => \N__17561\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__17567\,
            I => \N__17561\
        );

    \I__3945\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17557\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__17561\,
            I => \N__17554\
        );

    \I__3943\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17551\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__17557\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__17554\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17551\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17539\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17536\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__17542\,
            I => \N__17532\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17529\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17536\,
            I => \N__17526\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17523\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17520\
        );

    \I__3932\ : Span4Mux_h
    port map (
            O => \N__17529\,
            I => \N__17517\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__17526\,
            I => \N__17512\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17523\,
            I => \N__17512\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17520\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__17517\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__17512\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17500\
        );

    \I__3925\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17497\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__17503\,
            I => \N__17494\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17500\,
            I => \N__17490\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__17497\,
            I => \N__17487\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17484\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17481\
        );

    \I__3919\ : Span4Mux_h
    port map (
            O => \N__17490\,
            I => \N__17476\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__17487\,
            I => \N__17476\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__17484\,
            I => \N__17473\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__17481\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__17476\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__17473\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__3913\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17459\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17459\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__17464\,
            I => \N__17456\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__17459\,
            I => \N__17453\
        );

    \I__3909\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17449\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__17453\,
            I => \N__17446\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17443\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17449\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__17446\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17443\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__3903\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17432\
        );

    \I__3902\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17429\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17425\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__17429\,
            I => \N__17422\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17418\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__17425\,
            I => \N__17413\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__17422\,
            I => \N__17413\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17410\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17418\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__17413\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__17410\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__17403\,
            I => \N__17396\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17392\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \N__17388\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__17400\,
            I => \N__17384\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17367\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17367\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17367\
        );

    \I__3885\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17367\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17367\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17367\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17367\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17367\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17364\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__17364\,
            I => \N__17361\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__17361\,
            I => \Lab_UT.N_13_0\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17354\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17350\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17347\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \N__17344\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17350\,
            I => \N__17341\
        );

    \I__3872\ : Span4Mux_s0_v
    port map (
            O => \N__17347\,
            I => \N__17338\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17334\
        );

    \I__3870\ : Span4Mux_v
    port map (
            O => \N__17341\,
            I => \N__17329\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__17338\,
            I => \N__17329\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17326\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17334\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__17329\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17326\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17315\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17312\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__17315\,
            I => \N__17309\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17303\
        );

    \I__3860\ : Span12Mux_s5_v
    port map (
            O => \N__17309\,
            I => \N__17303\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17300\
        );

    \I__3858\ : Odrv12
    port map (
            O => \N__17303\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__17300\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17291\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17288\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17285\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17288\,
            I => \N__17279\
        );

    \I__3852\ : Span4Mux_v
    port map (
            O => \N__17285\,
            I => \N__17279\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17276\
        );

    \I__3850\ : Span4Mux_h
    port map (
            O => \N__17279\,
            I => \N__17273\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17270\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__17273\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__17270\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17260\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17257\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__17263\,
            I => \N__17254\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17260\,
            I => \N__17251\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17257\,
            I => \N__17248\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17245\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__17251\,
            I => \N__17242\
        );

    \I__3839\ : Span4Mux_h
    port map (
            O => \N__17248\,
            I => \N__17237\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17237\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__17242\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__17237\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__3835\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17228\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17225\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__17228\,
            I => \N__17220\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17225\,
            I => \N__17220\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__17220\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17211\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__17211\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17208\,
            I => \N__17198\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17198\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17206\,
            I => \N__17192\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17192\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17187\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17187\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17184\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17181\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__17192\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__17187\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__17184\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__17181\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17168\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17165\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17168\,
            I => \N__17162\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17159\
        );

    \I__3811\ : Span4Mux_h
    port map (
            O => \N__17162\,
            I => \N__17155\
        );

    \I__3810\ : Span4Mux_s2_v
    port map (
            O => \N__17159\,
            I => \N__17152\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17149\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__17155\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__17152\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__17149\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17139\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__17139\,
            I => \N__17136\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__17133\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_6\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__17130\,
            I => \N__17124\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17115\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17115\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17115\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17115\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17115\,
            I => \N__17112\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__17112\,
            I => \N__17109\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__17109\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__17106\,
            I => \N__17103\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17100\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17100\,
            I => \Lab_UT.didp.countrce3.q_5_3\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17091\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17091\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17091\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17084\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17080\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17084\,
            I => \N__17077\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17072\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17080\,
            I => \N__17069\
        );

    \I__3782\ : Span4Mux_s3_v
    port map (
            O => \N__17077\,
            I => \N__17066\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17061\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17075\,
            I => \N__17061\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__17072\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__17069\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__17066\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__17061\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17046\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17043\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17040\
        );

    \I__3772\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17036\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17046\,
            I => \N__17029\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17043\,
            I => \N__17029\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17029\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17024\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17036\,
            I => \N__17021\
        );

    \I__3766\ : Span4Mux_s3_v
    port map (
            O => \N__17029\,
            I => \N__17018\
        );

    \I__3765\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17013\
        );

    \I__3764\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17013\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17024\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__17021\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__17018\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17013\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16997\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16997\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16993\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16987\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__16996\,
            I => \N__16984\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__16993\,
            I => \N__16981\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16978\
        );

    \I__3752\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16973\
        );

    \I__3751\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16973\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__16987\,
            I => \N__16970\
        );

    \I__3749\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16967\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__16981\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__16978\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__16973\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__16970\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__16967\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3743\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16946\
        );

    \I__3742\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16946\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16946\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__16953\,
            I => \N__16943\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16938\
        );

    \I__3738\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16935\
        );

    \I__3737\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16932\
        );

    \I__3736\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16929\
        );

    \I__3735\ : Span4Mux_v
    port map (
            O => \N__16938\,
            I => \N__16926\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__16935\,
            I => \N__16923\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16920\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16917\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__16926\,
            I => \Lab_UT.LdMones\
        );

    \I__3730\ : Odrv12
    port map (
            O => \N__16923\,
            I => \Lab_UT.LdMones\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__16920\,
            I => \Lab_UT.LdMones\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__16917\,
            I => \Lab_UT.LdMones\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__16908\,
            I => \Lab_UT.didp.countrce3.un13_qPone_cascade_\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__16905\,
            I => \N__16901\
        );

    \I__3725\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16895\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16892\
        );

    \I__3723\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16889\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16899\,
            I => \N__16886\
        );

    \I__3721\ : InMux
    port map (
            O => \N__16898\,
            I => \N__16883\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__16895\,
            I => \N__16880\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__16892\,
            I => \N__16876\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16867\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N__16867\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__16883\,
            I => \N__16867\
        );

    \I__3715\ : Span4Mux_s3_v
    port map (
            O => \N__16880\,
            I => \N__16867\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16864\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__16876\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__16867\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__16864\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__16857\,
            I => \N__16854\
        );

    \I__3709\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16851\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__16851\,
            I => \Lab_UT.didp.countrce3.q_5_2\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__16848\,
            I => \N__16845\
        );

    \I__3706\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16835\
        );

    \I__3705\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16835\
        );

    \I__3704\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16835\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16832\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__16835\,
            I => \N__16829\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__16832\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__3700\ : Odrv12
    port map (
            O => \N__16829\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__3699\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16819\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16816\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \N__16812\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16809\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__16816\,
            I => \N__16806\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__16815\,
            I => \N__16803\
        );

    \I__3693\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16800\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__16809\,
            I => \N__16795\
        );

    \I__3691\ : Span4Mux_v
    port map (
            O => \N__16806\,
            I => \N__16795\
        );

    \I__3690\ : InMux
    port map (
            O => \N__16803\,
            I => \N__16792\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__16800\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__16795\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16792\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__3685\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16774\
        );

    \I__3684\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16769\
        );

    \I__3683\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16769\
        );

    \I__3682\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16766\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16761\
        );

    \I__3680\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16761\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__16774\,
            I => bu_rx_data_fast_1
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__16769\,
            I => bu_rx_data_fast_1
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__16766\,
            I => bu_rx_data_fast_1
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__16761\,
            I => bu_rx_data_fast_1
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__16752\,
            I => \N__16747\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \N__16742\
        );

    \I__3673\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16739\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16736\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__16746\,
            I => \N__16733\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16726\
        );

    \I__3669\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16726\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__16739\,
            I => \N__16721\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__16736\,
            I => \N__16721\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16717\
        );

    \I__3665\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16714\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__16731\,
            I => \N__16711\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16707\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__16721\,
            I => \N__16704\
        );

    \I__3661\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16701\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16696\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__16714\,
            I => \N__16696\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16691\
        );

    \I__3657\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16691\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__16707\,
            I => bu_rx_data_3_rep1
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__16704\,
            I => bu_rx_data_3_rep1
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__16701\,
            I => bu_rx_data_3_rep1
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__16696\,
            I => bu_rx_data_3_rep1
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__16691\,
            I => bu_rx_data_3_rep1
        );

    \I__3651\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16677\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__16674\,
            I => \Lab_UT.dictrl.g1_1Z0Z_1\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16668\,
            I => \N__16665\
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__16665\,
            I => \Lab_UT.dictrl.g2_1_0\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16659\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__16659\,
            I => \N__16656\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__16656\,
            I => \Lab_UT.dictrl.g2\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16646\
        );

    \I__3641\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16646\
        );

    \I__3640\ : InMux
    port map (
            O => \N__16651\,
            I => \N__16643\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16646\,
            I => \Lab_UT.didp.countrce3.ce_12_2_3\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__16643\,
            I => \Lab_UT.didp.countrce3.ce_12_2_3\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16635\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__16635\,
            I => \N__16631\
        );

    \I__3635\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16628\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__16631\,
            I => \N__16624\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__16628\,
            I => \N__16621\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__16627\,
            I => \N__16618\
        );

    \I__3631\ : Span4Mux_v
    port map (
            O => \N__16624\,
            I => \N__16613\
        );

    \I__3630\ : Span4Mux_s2_v
    port map (
            O => \N__16621\,
            I => \N__16613\
        );

    \I__3629\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16610\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__16613\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__16610\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__3626\ : CEMux
    port map (
            O => \N__16605\,
            I => \N__16601\
        );

    \I__3625\ : CEMux
    port map (
            O => \N__16604\,
            I => \N__16598\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__16601\,
            I => \N__16595\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__16598\,
            I => \N__16592\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__16595\,
            I => \N__16589\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__16592\,
            I => \N__16586\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__16589\,
            I => \N__16583\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__16586\,
            I => \N__16580\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__16583\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__16580\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__16575\,
            I => \Lab_UT.didp.un1_dicLdMones_0_cascade_\
        );

    \I__3615\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16569\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16566\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__16563\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__3611\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__16557\,
            I => \Lab_UT.dictrl.g0_2Z0Z_4\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__16554\,
            I => \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\
        );

    \I__3608\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16548\,
            I => \Lab_UT.dictrl.N_77_1_0\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__16545\,
            I => \Lab_UT.dictrl.N_77_1_0_cascade_\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16539\,
            I => \Lab_UT.dictrl.N_2353_0_0\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__16536\,
            I => \N__16528\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__16535\,
            I => \N__16525\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16520\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16520\
        );

    \I__3599\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16510\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16510\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16510\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16510\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__16520\,
            I => \N__16507\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__16519\,
            I => \N__16504\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__16510\,
            I => \N__16501\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__16507\,
            I => \N__16498\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16495\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__16501\,
            I => \N__16492\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__16498\,
            I => \buart__rx_shifter_fast_6\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__16495\,
            I => \buart__rx_shifter_fast_6\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__16492\,
            I => \buart__rx_shifter_fast_6\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__16485\,
            I => \N__16481\
        );

    \I__3585\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16470\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16470\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16470\
        );

    \I__3582\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16470\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16470\,
            I => \N__16466\
        );

    \I__3580\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16463\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__16466\,
            I => \N__16460\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__16463\,
            I => bu_rx_data_fast_7
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__16460\,
            I => bu_rx_data_fast_7
        );

    \I__3576\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16452\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__16452\,
            I => \Lab_UT.dictrl.state_fast_3\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16443\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16443\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16440\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__16440\,
            I => \Lab_UT.dictrl.g1_6\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__16437\,
            I => \Lab_UT.dictrl.m47_xZ0Z0_cascade_\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16429\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16424\
        );

    \I__3567\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16424\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16429\,
            I => \N__16417\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__16424\,
            I => \N__16417\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16412\
        );

    \I__3563\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16412\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__16417\,
            I => bu_rx_data_fast_4
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16412\,
            I => bu_rx_data_fast_4
        );

    \I__3560\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16401\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16401\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N__16398\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__16398\,
            I => \Lab_UT.dictrl.m30Z0Z_1\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16392\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__16392\,
            I => \Lab_UT.dictrl.N_81_0\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__16389\,
            I => \Lab_UT.dictrl.N_16_mux_0_cascade_\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16383\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__16383\,
            I => \Lab_UT.dictrl.N_113_0_0\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16373\
        );

    \I__3550\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16368\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16368\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16363\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16360\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16373\,
            I => \N__16356\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__16368\,
            I => \N__16353\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16350\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16347\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16363\,
            I => \N__16344\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16339\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16339\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__16356\,
            I => \N__16332\
        );

    \I__3538\ : Span4Mux_h
    port map (
            O => \N__16353\,
            I => \N__16332\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__16350\,
            I => \N__16332\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16347\,
            I => \N__16325\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__16344\,
            I => \N__16325\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__16339\,
            I => \N__16325\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__16332\,
            I => \N__16322\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__16325\,
            I => \Lab_UT.dictrl.state_2_rep1\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__16322\,
            I => \Lab_UT.dictrl.state_2_rep1\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__16317\,
            I => \Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16311\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16311\,
            I => \Lab_UT.dictrl.N_5_0\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16308\,
            I => \Lab_UT.dictrl.g2_2_cascade_\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16302\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16302\,
            I => \N__16298\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16295\
        );

    \I__3523\ : Odrv12
    port map (
            O => \N__16298\,
            I => \Lab_UT.dictrl.i9_mux_0\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16295\,
            I => \Lab_UT.dictrl.i9_mux_0\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16287\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__3519\ : Span4Mux_h
    port map (
            O => \N__16284\,
            I => \N__16280\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16277\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__16280\,
            I => \Lab_UT.dictrl.N_77_0\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__16277\,
            I => \Lab_UT.dictrl.N_77_0\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16267\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16264\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16261\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16267\,
            I => \N__16253\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__16264\,
            I => \N__16253\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16261\,
            I => \N__16250\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16247\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16242\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16242\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__16253\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__16250\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16247\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16242\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16230\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16230\,
            I => \Lab_UT.dictrl.g0_0Z0Z_1\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16224\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16224\,
            I => \N__16220\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16217\
        );

    \I__3497\ : Span12Mux_s6_h
    port map (
            O => \N__16220\,
            I => \N__16214\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16217\,
            I => \N__16211\
        );

    \I__3495\ : Odrv12
    port map (
            O => \N__16214\,
            I => \Lab_UT.dictrl.m30_0Z0Z_0\
        );

    \I__3494\ : Odrv12
    port map (
            O => \N__16211\,
            I => \Lab_UT.dictrl.m30_0Z0Z_0\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__16206\,
            I => \Lab_UT.dictrl.m25Z0Z_0_cascade_\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16200\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16200\,
            I => \N__16197\
        );

    \I__3490\ : Span4Mux_h
    port map (
            O => \N__16197\,
            I => \N__16194\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__16194\,
            I => \Lab_UT.dictrl.m59_ns_1_xZ0Z1\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__16191\,
            I => \Lab_UT.dictrl.N_81_1_cascade_\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16185\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__16185\,
            I => \Lab_UT.dictrl.N_113_1\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__16182\,
            I => \Lab_UT.dictrl.N_113_1_cascade_\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__3483\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16166\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16166\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16176\,
            I => \N__16166\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16173\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16166\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16156\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16153\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16150\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16145\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__16153\,
            I => \N__16145\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__16150\,
            I => \N__16142\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__16145\,
            I => \N__16139\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__16142\,
            I => \N__16136\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__16139\,
            I => \Lab_UT.dictrl.m59_ns_1\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__16136\,
            I => \Lab_UT.dictrl.m59_ns_1\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16128\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16125\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__16125\,
            I => \N__16122\
        );

    \I__3465\ : Odrv4
    port map (
            O => \N__16122\,
            I => \Lab_UT.dictrl.state_fast_2\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__16119\,
            I => \N__16116\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16107\
        );

    \I__3462\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16107\
        );

    \I__3461\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16107\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16107\,
            I => \N__16103\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16100\
        );

    \I__3458\ : Span4Mux_h
    port map (
            O => \N__16103\,
            I => \N__16097\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__16100\,
            I => \N__16094\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__16097\,
            I => \N__16091\
        );

    \I__3455\ : Sp12to4
    port map (
            O => \N__16094\,
            I => \N__16088\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__16091\,
            I => \Lab_UT.dictrl.g0_17_0\
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__16088\,
            I => \Lab_UT.dictrl.g0_17_0\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16074\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16074\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16074\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__16074\,
            I => \N__16070\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16067\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__16070\,
            I => \N__16064\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16067\,
            I => \N__16061\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__16064\,
            I => \N__16057\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__16061\,
            I => \N__16054\
        );

    \I__3443\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16051\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__16057\,
            I => \Lab_UT.dictrl.g0_17_1\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__16054\,
            I => \Lab_UT.dictrl.g0_17_1\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__16051\,
            I => \Lab_UT.dictrl.g0_17_1\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16040\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16036\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__16040\,
            I => \N__16031\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16027\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16024\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16021\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16018\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__16031\,
            I => \N__16015\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16012\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__16027\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__16024\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__16021\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__16018\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__16015\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16012\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3424\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15995\
        );

    \I__3423\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15990\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__15995\,
            I => \N__15987\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15983\
        );

    \I__3420\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15980\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15977\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__15987\,
            I => \N__15974\
        );

    \I__3417\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15971\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__15983\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__15980\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__15977\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__15974\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__15971\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3411\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15942\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15942\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15942\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15942\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15942\
        );

    \I__3406\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15942\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__15942\,
            I => \N__15938\
        );

    \I__3404\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15935\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__15938\,
            I => \N__15932\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__15935\,
            I => \Lab_UT.didp.un18_ce\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__15932\,
            I => \Lab_UT.didp.un18_ce\
        );

    \I__3400\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15924\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__15924\,
            I => \N__15921\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__15921\,
            I => \Lab_UT.LdSones_i_3\
        );

    \I__3397\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15914\
        );

    \I__3396\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15911\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15908\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__15911\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__15908\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__15903\,
            I => \N__15898\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__15902\,
            I => \N__15894\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15887\
        );

    \I__3389\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15887\
        );

    \I__3388\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15887\
        );

    \I__3387\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15884\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__15887\,
            I => \N__15881\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15878\
        );

    \I__3384\ : Odrv12
    port map (
            O => \N__15881\,
            I => \Lab_UT.LdStens\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__15878\,
            I => \Lab_UT.LdStens\
        );

    \I__3382\ : CEMux
    port map (
            O => \N__15873\,
            I => \N__15858\
        );

    \I__3381\ : CEMux
    port map (
            O => \N__15872\,
            I => \N__15858\
        );

    \I__3380\ : CEMux
    port map (
            O => \N__15871\,
            I => \N__15858\
        );

    \I__3379\ : CEMux
    port map (
            O => \N__15870\,
            I => \N__15858\
        );

    \I__3378\ : CEMux
    port map (
            O => \N__15869\,
            I => \N__15858\
        );

    \I__3377\ : GlobalMux
    port map (
            O => \N__15858\,
            I => \N__15855\
        );

    \I__3376\ : gio2CtrlBuf
    port map (
            O => \N__15855\,
            I => bu_rx_data_rdy_0_g
        );

    \I__3375\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15849\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__15849\,
            I => \Lab_UT.didp.countrce1.un13_qPone\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__15846\,
            I => \Lab_UT.didp.countrce1.q_5_2_cascade_\
        );

    \I__3372\ : InMux
    port map (
            O => \N__15843\,
            I => \N__15839\
        );

    \I__3371\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15836\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__15839\,
            I => \N__15833\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15828\
        );

    \I__3368\ : Span4Mux_v
    port map (
            O => \N__15833\,
            I => \N__15825\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15820\
        );

    \I__3366\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15820\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__15828\,
            I => \N__15817\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__15825\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15820\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__15817\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__3361\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15807\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__15807\,
            I => \N__15803\
        );

    \I__3359\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15798\
        );

    \I__3358\ : Span4Mux_v
    port map (
            O => \N__15803\,
            I => \N__15795\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15790\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15790\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15798\,
            I => \N__15787\
        );

    \I__3354\ : Span4Mux_s1_v
    port map (
            O => \N__15795\,
            I => \N__15784\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__15790\,
            I => \N__15779\
        );

    \I__3352\ : Sp12to4
    port map (
            O => \N__15787\,
            I => \N__15779\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__15784\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3350\ : Odrv12
    port map (
            O => \N__15779\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3349\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15771\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__15771\,
            I => \N__15768\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__15768\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15762\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__15762\,
            I => \Lab_UT.un1_idle_5_0_iclkZ0\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__15759\,
            I => \N__15756\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15753\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__15753\,
            I => \N__15748\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15745\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15741\
        );

    \I__3339\ : Span4Mux_v
    port map (
            O => \N__15748\,
            I => \N__15736\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15736\
        );

    \I__3337\ : SRMux
    port map (
            O => \N__15744\,
            I => \N__15733\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__15741\,
            I => \N__15730\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__15736\,
            I => \N__15724\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__15733\,
            I => \N__15724\
        );

    \I__3333\ : Span12Mux_v
    port map (
            O => \N__15730\,
            I => \N__15721\
        );

    \I__3332\ : IoInMux
    port map (
            O => \N__15729\,
            I => \N__15718\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__15724\,
            I => \N__15715\
        );

    \I__3330\ : Odrv12
    port map (
            O => \N__15721\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__15718\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__15715\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__15708\,
            I => \Lab_UT.un1_armed_2_0_iso_iZ0_cascade_\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15701\
        );

    \I__3325\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15698\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__15701\,
            I => \G_192\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__15698\,
            I => \G_192\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__15693\,
            I => \Lab_UT.dictrl.N_113_cascade_\
        );

    \I__3321\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__3319\ : Span4Mux_h
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__15681\,
            I => \Lab_UT.didp.did_alarmMatch_7\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__15678\,
            I => \Lab_UT.didp.did_alarmMatch_4_cascade_\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15672\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__15672\,
            I => \Lab_UT.didp.did_alarmMatch_5\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__15669\,
            I => \Lab_UT.did_alarmMatch_13_cascade_\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__15666\,
            I => \Lab_UT.dictrl.alarmstate_1_0_cascade_\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15660\,
            I => \Lab_UT.did_alarmMatch_13\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__15657\,
            I => \G_183_cascade_\
        );

    \I__3309\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15648\
        );

    \I__3308\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15648\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__15648\,
            I => \N__15645\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__15645\,
            I => \Lab_UT.did_alarmMatch_12\
        );

    \I__3305\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15639\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__15639\,
            I => \N__15636\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__15636\,
            I => \Lab_UT.didp.countrce2.un13_qPone\
        );

    \I__3302\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15628\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15622\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15622\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__15628\,
            I => \N__15619\
        );

    \I__3298\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15614\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15611\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__15619\,
            I => \N__15608\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15603\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15603\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15614\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__15611\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__15608\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__15603\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15591\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15591\,
            I => \N__15588\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__15588\,
            I => \Lab_UT.didp.countrce2.q_5_2\
        );

    \I__3286\ : IoInMux
    port map (
            O => \N__15585\,
            I => \N__15579\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15575\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15571\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15568\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15579\,
            I => \N__15565\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15562\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__15575\,
            I => \N__15559\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15556\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__15571\,
            I => \N__15553\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15568\,
            I => \N__15550\
        );

    \I__3276\ : Span4Mux_s0_h
    port map (
            O => \N__15565\,
            I => \N__15547\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15562\,
            I => \N__15544\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__15559\,
            I => \N__15541\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__15556\,
            I => \N__15538\
        );

    \I__3272\ : Span4Mux_v
    port map (
            O => \N__15553\,
            I => \N__15533\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__15550\,
            I => \N__15533\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__15547\,
            I => \N__15530\
        );

    \I__3269\ : Span4Mux_v
    port map (
            O => \N__15544\,
            I => \N__15527\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__15541\,
            I => rst
        );

    \I__3267\ : Odrv12
    port map (
            O => \N__15538\,
            I => rst
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__15533\,
            I => rst
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15530\,
            I => rst
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__15527\,
            I => rst
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15509\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15506\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15509\,
            I => \G_184\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15506\,
            I => \G_184\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__15501\,
            I => \N__15497\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15494\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15490\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15494\,
            I => \N__15487\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15484\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15490\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__15487\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15484\,
            I => \Lab_UT.alarmstate_0_sqmuxa_1\
        );

    \I__3250\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15473\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15470\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__15473\,
            I => \N__15462\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15470\,
            I => \N__15462\
        );

    \I__3246\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15455\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15455\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15455\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__15462\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__15455\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15447\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15447\,
            I => \Lab_UT.didp.countrce2.q_5_3\
        );

    \I__3239\ : InMux
    port map (
            O => \N__15444\,
            I => \N__15441\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__15438\,
            I => \Lab_UT.didp.countrce2.q_5_0\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__15435\,
            I => \N__15427\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15434\,
            I => \N__15423\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15414\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15414\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15414\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15414\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15427\,
            I => \N__15408\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15408\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15405\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15414\,
            I => \N__15402\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15399\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15408\,
            I => \N__15396\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15405\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__15402\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15399\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__15396\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__15387\,
            I => \N__15382\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15375\
        );

    \I__3218\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15372\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15369\
        );

    \I__3216\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15364\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15364\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15359\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15359\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__15375\,
            I => \N__15356\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15372\,
            I => \N__15353\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15369\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__15364\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__15359\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3207\ : Odrv12
    port map (
            O => \N__15356\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__15353\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15335\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15332\
        );

    \I__3203\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15329\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15326\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15323\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15335\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15332\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__15329\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__15326\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__15323\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15309\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15309\,
            I => \Lab_UT.didp.regrce3.did_alarmMatch_3\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15303\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15303\,
            I => \Lab_UT.didp.did_alarmMatch_0\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__15300\,
            I => \Lab_UT.didp.did_alarmMatch_1_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15294\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__15294\,
            I => \N__15291\
        );

    \I__3188\ : Odrv4
    port map (
            O => \N__15291\,
            I => \Lab_UT.didp.did_alarmMatch_2\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__15288\,
            I => \N__15283\
        );

    \I__3186\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15277\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15277\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15272\
        );

    \I__3183\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15272\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15267\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15267\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__15267\,
            I => \N__15264\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__15264\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15261\,
            I => \N__15256\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__15260\,
            I => \N__15253\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15247\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15247\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15242\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15242\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__15247\,
            I => \N__15239\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15236\
        );

    \I__3170\ : Span4Mux_h
    port map (
            O => \N__15239\,
            I => \N__15233\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__15236\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__15233\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__15228\,
            I => \N__15223\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__15227\,
            I => \N__15220\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__15226\,
            I => \N__15215\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15208\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15208\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15208\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15203\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15203\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15208\,
            I => \Lab_UT.didp.un24_ce_2\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__15203\,
            I => \Lab_UT.didp.un24_ce_2\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15193\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15190\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__15196\,
            I => \N__15185\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15179\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15190\,
            I => \N__15179\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15176\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15171\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15171\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15168\
        );

    \I__3148\ : Span4Mux_s2_v
    port map (
            O => \N__15179\,
            I => \N__15163\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15176\,
            I => \N__15163\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15171\,
            I => \N__15158\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15158\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__15163\,
            I => \Lab_UT.LdMtens\
        );

    \I__3143\ : Odrv12
    port map (
            O => \N__15158\,
            I => \Lab_UT.LdMtens\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__15153\,
            I => \N__15150\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15147\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15147\,
            I => \N__15144\
        );

    \I__3139\ : Span4Mux_h
    port map (
            O => \N__15144\,
            I => \N__15141\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__15141\,
            I => \Lab_UT.didp.countrce4.un20_qPone\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15133\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15130\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15127\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15133\,
            I => \N__15124\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15130\,
            I => \N__15119\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15127\,
            I => \N__15119\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__15124\,
            I => \N__15113\
        );

    \I__3130\ : Span4Mux_v
    port map (
            O => \N__15119\,
            I => \N__15113\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15110\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__15113\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15110\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__15105\,
            I => \Lab_UT.didp.countrce4.q_5_3_cascade_\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15099\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15099\,
            I => \N__15094\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15089\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15089\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__15094\,
            I => \N__15086\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__15089\,
            I => \N__15083\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__15086\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__15083\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15075\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__15075\,
            I => \Lab_UT.didp.countrce2.q_5_1\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__15072\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15066\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15066\,
            I => \Lab_UT.didp.reset_12_1_3\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15057\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15052\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15052\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15047\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15044\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15052\,
            I => \N__15041\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15036\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15036\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15047\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__15044\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__3102\ : Odrv12
    port map (
            O => \N__15041\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15036\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__15027\,
            I => \Lab_UT.didp.ce_12_3_cascade_\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__15024\,
            I => \N__15021\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15006\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15006\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15019\,
            I => \N__14992\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14992\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15017\,
            I => \N__14992\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15016\,
            I => \N__14992\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15015\,
            I => \N__14992\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15014\,
            I => \N__14992\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15013\,
            I => \N__14989\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15012\,
            I => \N__14986\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14983\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15006\,
            I => \N__14980\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15005\,
            I => \N__14977\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14972\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14972\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__14986\,
            I => \N__14969\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__14983\,
            I => \N__14966\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__14980\,
            I => \N__14960\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__14977\,
            I => \N__14960\
        );

    \I__3079\ : Span4Mux_s2_v
    port map (
            O => \N__14972\,
            I => \N__14957\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__14969\,
            I => \N__14952\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__14966\,
            I => \N__14952\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14949\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__14960\,
            I => \N__14944\
        );

    \I__3074\ : Span4Mux_h
    port map (
            O => \N__14957\,
            I => \N__14944\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__14952\,
            I => \oneSecStrb\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__14949\,
            I => \oneSecStrb\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__14944\,
            I => \oneSecStrb\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__14937\,
            I => \Lab_UT.didp.countrce2.un20_qPone_cascade_\
        );

    \I__3069\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14931\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__14931\,
            I => \Lab_UT.didp.countrce4.q_5_0\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__14928\,
            I => \N__14925\
        );

    \I__3066\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14921\
        );

    \I__3065\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14918\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__14921\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__14918\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__14913\,
            I => \Lab_UT.dictrl.g0_17_0_cascade_\
        );

    \I__3061\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14907\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__14907\,
            I => \N__14904\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__14904\,
            I => \Lab_UT.dictrl.g2_0_0\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__14901\,
            I => \N__14897\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14891\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14891\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14888\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14883\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14883\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__14883\,
            I => bu_rx_data_fast_3
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__14880\,
            I => \Lab_UT.dictrl.g0_2Z0Z_5_cascade_\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14877\,
            I => \N__14874\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14874\,
            I => \N__14871\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__14871\,
            I => \Lab_UT.dictrl.g2_0\
        );

    \I__3047\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14865\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__14865\,
            I => \Lab_UT.dictrl.g1_1\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__14862\,
            I => \Lab_UT.dictrl.g2_0_cascade_\
        );

    \I__3044\ : InMux
    port map (
            O => \N__14859\,
            I => \N__14856\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14856\,
            I => \Lab_UT.dictrl.N_90_0_0_0\
        );

    \I__3042\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__14850\,
            I => \Lab_UT.dictrl.m40_N_5_mux_0\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__14847\,
            I => \Lab_UT.dictrl.g2Z0Z_1_cascade_\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14841\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__14841\,
            I => \N__14838\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__14838\,
            I => \N__14834\
        );

    \I__3036\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14831\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__14834\,
            I => \Lab_UT.dictrl.g1_0\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__14831\,
            I => \Lab_UT.dictrl.g1_0\
        );

    \I__3033\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14823\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__14823\,
            I => \Lab_UT.dictrl.g0_17_a6_2_1\
        );

    \I__3031\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14817\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14817\,
            I => \N__14814\
        );

    \I__3029\ : Odrv12
    port map (
            O => \N__14814\,
            I => \Lab_UT.dictrl.g0_17_a6_3_6\
        );

    \I__3028\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__14808\,
            I => \Lab_UT.dictrl.g0_17_a6_3_8\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__14805\,
            I => \Lab_UT.dictrl.N_22_cascade_\
        );

    \I__3025\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14790\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14790\
        );

    \I__3023\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14790\
        );

    \I__3022\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14790\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14787\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__14787\,
            I => \Lab_UT.dictrl.N_90_0\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__14784\,
            I => \N__14778\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__14783\,
            I => \N__14775\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__14782\,
            I => \N__14772\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__14781\,
            I => \N__14769\
        );

    \I__3015\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14764\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14764\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14772\,
            I => \N__14759\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14759\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14754\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__14759\,
            I => \N__14754\
        );

    \I__3009\ : Odrv12
    port map (
            O => \N__14754\,
            I => \Lab_UT.dictrl.N_95_0\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__14751\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14745\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__14745\,
            I => \N__14742\
        );

    \I__3005\ : Odrv12
    port map (
            O => \N__14742\,
            I => \Lab_UT.LdStens_i_3\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__14739\,
            I => \N__14735\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \N__14731\
        );

    \I__3002\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14728\
        );

    \I__3001\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14725\
        );

    \I__3000\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14722\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__14728\,
            I => \N__14717\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__14725\,
            I => \N__14717\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14722\,
            I => \Lab_UT.dictrl.state_fast_1\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__14717\,
            I => \Lab_UT.dictrl.state_fast_1\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__14712\,
            I => \Lab_UT.dictrl.N_95_0_0_cascade_\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__14709\,
            I => \Lab_UT.dictrl.g0_3_0_cascade_\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__14706\,
            I => \Lab_UT.dictrl.g4_cascade_\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__14703\,
            I => \Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14697\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__14697\,
            I => \Lab_UT.dictrl.g2_5\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14688\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14681\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14681\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14681\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14688\,
            I => \N__14678\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__14681\,
            I => \Lab_UT.dicRun_2\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__14678\,
            I => \Lab_UT.dicRun_2\
        );

    \I__2982\ : InMux
    port map (
            O => \N__14673\,
            I => \N__14670\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14670\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__2980\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14664\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__14664\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14655\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14655\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14655\,
            I => \N__14650\
        );

    \I__2975\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14647\
        );

    \I__2974\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14644\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__14650\,
            I => \N__14641\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14647\,
            I => \N__14636\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__14644\,
            I => \N__14636\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__14641\,
            I => \N__14633\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__14636\,
            I => \N__14630\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__14633\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__14630\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14622\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__14622\,
            I => \Lab_UT.un1_idle_1_0_iclkZ0\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__14619\,
            I => \G_186_cascade_\
        );

    \I__2963\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14611\
        );

    \I__2962\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14606\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14606\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14611\,
            I => \G_191\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__14606\,
            I => \G_191\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__14601\,
            I => \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_\
        );

    \I__2957\ : InMux
    port map (
            O => \N__14598\,
            I => \N__14595\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__14595\,
            I => \N__14592\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__14592\,
            I => \Lab_UT.dictrl.G_10_1\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__14589\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__14586\,
            I => \Lab_UT.dictrl.N_21_0_cascade_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14573\
        );

    \I__2951\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14573\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14573\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14558\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14555\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14548\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14548\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14548\
        );

    \I__2944\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14539\
        );

    \I__2943\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14539\
        );

    \I__2942\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14539\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14539\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14536\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14531\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14531\
        );

    \I__2937\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14526\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14526\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__14558\,
            I => \N__14521\
        );

    \I__2934\ : Span4Mux_s1_v
    port map (
            O => \N__14555\,
            I => \N__14521\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14548\,
            I => \N__14518\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14515\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14536\,
            I => \Lab_UT.i16_mux\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14531\,
            I => \Lab_UT.i16_mux\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14526\,
            I => \Lab_UT.i16_mux\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__14521\,
            I => \Lab_UT.i16_mux\
        );

    \I__2927\ : Odrv12
    port map (
            O => \N__14518\,
            I => \Lab_UT.i16_mux\
        );

    \I__2926\ : Odrv12
    port map (
            O => \N__14515\,
            I => \Lab_UT.i16_mux\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14499\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14499\,
            I => \Lab_UT.dictrl.i18_mux\
        );

    \I__2923\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14493\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14493\,
            I => \Lab_UT.dispString.dOut_RNO_1Z0Z_1\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__14490\,
            I => \N__14484\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__14489\,
            I => \N__14477\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__14488\,
            I => \N__14473\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14466\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14466\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14459\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14459\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14459\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14450\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14447\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14442\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14442\
        );

    \I__2909\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14436\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14436\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14466\,
            I => \N__14433\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14430\
        );

    \I__2905\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14425\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14425\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14422\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14415\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14415\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14415\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14408\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14447\,
            I => \N__14408\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14408\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14404\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__14436\,
            I => \N__14399\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__14433\,
            I => \N__14399\
        );

    \I__2893\ : Span4Mux_h
    port map (
            O => \N__14430\,
            I => \N__14394\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14425\,
            I => \N__14394\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14422\,
            I => \N__14391\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14415\,
            I => \N__14386\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__14408\,
            I => \N__14386\
        );

    \I__2888\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14383\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__14404\,
            I => \N__14376\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__14399\,
            I => \N__14376\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__14394\,
            I => \N__14376\
        );

    \I__2884\ : Odrv12
    port map (
            O => \N__14391\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__14386\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14383\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__14376\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14358\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__14366\,
            I => \N__14353\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14350\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__14364\,
            I => \N__14347\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__14363\,
            I => \N__14344\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14341\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__14361\,
            I => \N__14337\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14358\,
            I => \N__14331\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14324\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14324\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14324\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__14350\,
            I => \N__14321\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14316\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14316\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14341\,
            I => \N__14313\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14303\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14337\,
            I => \N__14303\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14303\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14298\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14298\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__14331\,
            I => \N__14292\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14324\,
            I => \N__14292\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__14321\,
            I => \N__14287\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14316\,
            I => \N__14287\
        );

    \I__2856\ : Span4Mux_h
    port map (
            O => \N__14313\,
            I => \N__14284\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14277\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14277\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14277\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14303\,
            I => \N__14272\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14272\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14269\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__14292\,
            I => \N__14264\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__14287\,
            I => \N__14264\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__14284\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14277\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__14272\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14269\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__14264\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14250\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14247\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__14247\,
            I => \N__14244\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__14244\,
            I => \Lab_UT.dispString.m49_ns_1\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__14241\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__14238\,
            I => \Lab_UT.didp.countrce1.q_5_3_cascade_\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__14235\,
            I => \N__14226\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__14234\,
            I => \N__14223\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14220\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__14232\,
            I => \N__14217\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__14231\,
            I => \N__14214\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__14230\,
            I => \N__14211\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__14229\,
            I => \N__14208\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14199\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14199\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14199\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14199\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14196\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14191\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14191\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14199\,
            I => \Lab_UT.sec1_3\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14196\,
            I => \Lab_UT.sec1_3\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14191\,
            I => \Lab_UT.sec1_3\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14181\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__14181\,
            I => \N__14176\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14173\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14170\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__14176\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14173\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14170\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14163\,
            I => \N__14160\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14160\,
            I => \N__14156\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14152\
        );

    \I__2809\ : Span4Mux_s0_v
    port map (
            O => \N__14156\,
            I => \N__14149\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14155\,
            I => \N__14146\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14152\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__14149\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14146\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14139\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14129\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14126\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14134\,
            I => \N__14121\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14133\,
            I => \N__14116\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14116\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14129\,
            I => \N__14111\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14126\,
            I => \N__14111\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14108\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14103\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14103\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14116\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__14111\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14108\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__14103\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__14094\,
            I => \Lab_UT.didp.countrce4.un13_qPone_cascade_\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__14091\,
            I => \Lab_UT.didp.countrce4.q_5_2_cascade_\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__14088\,
            I => \Lab_UT.dictrl.N_95_cascade_\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14081\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14078\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14073\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14070\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14067\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14076\,
            I => \N__14064\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__14073\,
            I => \N__14052\
        );

    \I__2779\ : Span4Mux_s2_h
    port map (
            O => \N__14070\,
            I => \N__14052\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14067\,
            I => \N__14052\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__14064\,
            I => \N__14049\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14038\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14038\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14038\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14038\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14038\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__14052\,
            I => \uu2.N_101\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__14049\,
            I => \uu2.N_101\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14038\,
            I => \uu2.N_101\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__14031\,
            I => \N__14027\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14030\,
            I => \N__14024\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14020\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14015\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14015\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__14020\,
            I => \N__14012\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14015\,
            I => \N__14009\
        );

    \I__2761\ : Span4Mux_s2_v
    port map (
            O => \N__14012\,
            I => \N__14006\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__14009\,
            I => \N__14003\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__14006\,
            I => \uu2.N_111\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__14003\,
            I => \uu2.N_111\
        );

    \I__2757\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13994\
        );

    \I__2756\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13991\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__13994\,
            I => \N__13987\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__13991\,
            I => \N__13984\
        );

    \I__2753\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13981\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__13987\,
            I => \N__13977\
        );

    \I__2751\ : Span4Mux_s1_h
    port map (
            O => \N__13984\,
            I => \N__13972\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__13981\,
            I => \N__13972\
        );

    \I__2749\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13969\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__13977\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__13972\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__13969\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__13962\,
            I => \N__13959\
        );

    \I__2744\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13956\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13950\
        );

    \I__2742\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13945\
        );

    \I__2741\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13945\
        );

    \I__2740\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13942\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__13950\,
            I => \N__13937\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13937\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__13942\,
            I => \N__13932\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__13937\,
            I => \N__13932\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__13932\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2734\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13925\
        );

    \I__2733\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13922\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__13925\,
            I => \N__13919\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13912\
        );

    \I__2730\ : Span4Mux_s3_v
    port map (
            O => \N__13919\,
            I => \N__13909\
        );

    \I__2729\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13906\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13901\
        );

    \I__2727\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13901\
        );

    \I__2726\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13898\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__13912\,
            I => \N__13893\
        );

    \I__2724\ : Span4Mux_h
    port map (
            O => \N__13909\,
            I => \N__13893\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__13906\,
            I => \N__13888\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__13901\,
            I => \N__13888\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__13898\,
            I => \o_One_Sec_Pulse\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__13893\,
            I => \o_One_Sec_Pulse\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__13888\,
            I => \o_One_Sec_Pulse\
        );

    \I__2718\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13878\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13878\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__2716\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13872\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__13872\,
            I => \N__13868\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13865\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__13868\,
            I => \N__13862\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__13865\,
            I => \N__13857\
        );

    \I__2711\ : Span4Mux_v
    port map (
            O => \N__13862\,
            I => \N__13854\
        );

    \I__2710\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13849\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13849\
        );

    \I__2708\ : Span12Mux_s9_v
    port map (
            O => \N__13857\,
            I => \N__13846\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__13854\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13849\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2705\ : Odrv12
    port map (
            O => \N__13846\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13836\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__13836\,
            I => \N__13832\
        );

    \I__2702\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13829\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__13832\,
            I => \N__13826\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__13829\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__13826\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2698\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13818\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__13818\,
            I => \N__13815\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__13815\,
            I => \N__13812\
        );

    \I__2695\ : Span4Mux_s2_v
    port map (
            O => \N__13812\,
            I => \N__13809\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__13809\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__2693\ : InMux
    port map (
            O => \N__13806\,
            I => \N__13803\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__13803\,
            I => \N__13800\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__13800\,
            I => \N__13797\
        );

    \I__2690\ : Span4Mux_s2_v
    port map (
            O => \N__13797\,
            I => \N__13794\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__13794\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__13791\,
            I => \N__13788\
        );

    \I__2687\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13785\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13782\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__13782\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2684\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13766\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13766\
        );

    \I__2682\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13766\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13757\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13757\
        );

    \I__2679\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13757\
        );

    \I__2678\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13757\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13766\,
            I => \Lab_UT.sec1_2\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__13757\,
            I => \Lab_UT.sec1_2\
        );

    \I__2675\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13738\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13738\
        );

    \I__2672\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13729\
        );

    \I__2671\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13729\
        );

    \I__2670\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13729\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13729\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__13743\,
            I => \Lab_UT.sec1_1\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13738\,
            I => \Lab_UT.sec1_1\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13729\,
            I => \Lab_UT.sec1_1\
        );

    \I__2665\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13709\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13709\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13709\
        );

    \I__2662\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13700\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13700\
        );

    \I__2660\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13700\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13700\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__13709\,
            I => \N__13697\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__13700\,
            I => \N__13694\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__13697\,
            I => \Lab_UT.sec1_0\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__13694\,
            I => \Lab_UT.sec1_0\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13686\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13686\,
            I => \N__13683\
        );

    \I__2652\ : Odrv12
    port map (
            O => \N__13683\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__13680\,
            I => \N__13675\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__13679\,
            I => \N__13672\
        );

    \I__2649\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13659\
        );

    \I__2648\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13659\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13659\
        );

    \I__2646\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13659\
        );

    \I__2645\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13659\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__13659\,
            I => \N__13655\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__13658\,
            I => \N__13651\
        );

    \I__2642\ : Span4Mux_s0_v
    port map (
            O => \N__13655\,
            I => \N__13648\
        );

    \I__2641\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13643\
        );

    \I__2640\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13643\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__13648\,
            I => \Lab_UT.min1_2\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__13643\,
            I => \Lab_UT.min1_2\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13623\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13623\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13623\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13623\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13623\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13618\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13622\,
            I => \N__13613\
        );

    \I__2630\ : InMux
    port map (
            O => \N__13621\,
            I => \N__13613\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__13618\,
            I => \Lab_UT.min1_0\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__13613\,
            I => \Lab_UT.min1_0\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__13608\,
            I => \N__13604\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13592\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13592\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13592\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13583\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13583\
        );

    \I__2621\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13583\
        );

    \I__2620\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13583\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13592\,
            I => \Lab_UT.min2_1\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__13583\,
            I => \Lab_UT.min2_1\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13565\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13565\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13576\,
            I => \N__13565\
        );

    \I__2614\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13556\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13556\
        );

    \I__2612\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13556\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13556\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__13565\,
            I => \Lab_UT.min2_0\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13556\,
            I => \Lab_UT.min2_0\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__13551\,
            I => \N__13544\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__13550\,
            I => \N__13541\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__13549\,
            I => \N__13538\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__13548\,
            I => \N__13534\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__13547\,
            I => \N__13531\
        );

    \I__2603\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13521\
        );

    \I__2602\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13521\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13521\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13521\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13514\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13514\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13514\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13521\,
            I => \Lab_UT.min2_2\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__13514\,
            I => \Lab_UT.min2_2\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__13509\,
            I => \Lab_UT.dispString.N_18_0_cascade_\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13503\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__13503\,
            I => \N__13500\
        );

    \I__2591\ : Span4Mux_v
    port map (
            O => \N__13500\,
            I => \N__13497\
        );

    \I__2590\ : Span4Mux_h
    port map (
            O => \N__13497\,
            I => \N__13494\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__13494\,
            I => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13488\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13488\,
            I => \Lab_UT.dictrl.g0_17_a6_1_7\
        );

    \I__2586\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13482\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__13482\,
            I => \Lab_UT.dictrl.g0_17_a6_1Z0Z_6\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__13479\,
            I => \Lab_UT.dictrl.g0_17_a6_1_5_cascade_\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__13476\,
            I => \Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13473\,
            I => \N__13470\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__13470\,
            I => \Lab_UT.dictrl.g0_17_a6_2\
        );

    \I__2580\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13464\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13464\,
            I => \Lab_UT.dictrl.N_19\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13461\,
            I => \N__13458\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__13458\,
            I => \Lab_UT.dictrl.g0_17_o6_1Z0Z_5\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__13455\,
            I => \N__13449\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13440\
        );

    \I__2574\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13440\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13440\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13440\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13440\,
            I => \N__13434\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13427\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13427\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13437\,
            I => \N__13427\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__13434\,
            I => \Lab_UT.min2_3\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13427\,
            I => \Lab_UT.min2_3\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__13422\,
            I => \N__13416\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__13421\,
            I => \N__13411\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__13420\,
            I => \N__13408\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__13419\,
            I => \N__13405\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13393\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13393\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13393\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13393\
        );

    \I__2557\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13393\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13388\
        );

    \I__2555\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13388\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13393\,
            I => \N__13385\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13388\,
            I => \N__13382\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__13385\,
            I => \Lab_UT.min1_3\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__13382\,
            I => \Lab_UT.min1_3\
        );

    \I__2550\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13374\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13374\,
            I => \Lab_UT.dictrl.g1Z0Z_5\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13371\,
            I => \Lab_UT.dictrl.g1_cascade_\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__13368\,
            I => \Lab_UT.dictrl.g0_2_3_cascade_\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13361\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13358\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13361\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13358\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13353\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13350\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13347\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13344\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13331\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13331\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13331\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13328\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13331\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13328\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13323\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13311\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13311\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13311\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2526\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13299\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13299\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13299\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__13296\,
            I => \N__13292\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13295\,
            I => \N__13289\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13286\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13289\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13286\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13275\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13275\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13275\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13269\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__13269\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13263\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13263\,
            I => \N__13260\
        );

    \I__2511\ : Span4Mux_s2_h
    port map (
            O => \N__13260\,
            I => \N__13257\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__13257\,
            I => \N__13252\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13249\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13246\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__13252\,
            I => \L3_tx_data_1\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13249\,
            I => \L3_tx_data_1\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13246\,
            I => \L3_tx_data_1\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13236\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13236\,
            I => \Lab_UT.dispString.m42_ns_1\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__13230\,
            I => \N__13227\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__13227\,
            I => vbuf_tx_data_6
        );

    \I__2499\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__13221\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__13218\,
            I => \N__13213\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13207\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13207\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13202\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13202\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13207\,
            I => \N__13194\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13202\,
            I => \N__13194\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13189\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13189\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13199\,
            I => \N__13177\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__13194\,
            I => \N__13172\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13189\,
            I => \N__13172\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13155\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13187\,
            I => \N__13155\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13186\,
            I => \N__13155\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13155\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13155\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13155\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13155\
        );

    \I__2478\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13155\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13152\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13149\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__13172\,
            I => \N__13146\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13155\,
            I => \N__13141\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__13152\,
            I => \N__13141\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13149\,
            I => vbuf_tx_data_rdy
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__13146\,
            I => vbuf_tx_data_rdy
        );

    \I__2470\ : Odrv12
    port map (
            O => \N__13141\,
            I => vbuf_tx_data_rdy
        );

    \I__2469\ : InMux
    port map (
            O => \N__13134\,
            I => \N__13131\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__13128\,
            I => vbuf_tx_data_7
        );

    \I__2466\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13122\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13122\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__2464\ : CEMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13116\,
            I => \N__13112\
        );

    \I__2462\ : CEMux
    port map (
            O => \N__13115\,
            I => \N__13109\
        );

    \I__2461\ : Span4Mux_v
    port map (
            O => \N__13112\,
            I => \N__13106\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13109\,
            I => \N__13103\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__13106\,
            I => \N__13100\
        );

    \I__2458\ : Span4Mux_v
    port map (
            O => \N__13103\,
            I => \N__13097\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__13100\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__13097\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__13091\,
            I => \N__13081\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13075\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13070\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13070\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__13085\,
            I => \N__13065\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13056\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13056\
        );

    \I__2447\ : InMux
    port map (
            O => \N__13080\,
            I => \N__13056\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13079\,
            I => \N__13056\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__13078\,
            I => \N__13052\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13075\,
            I => \N__13049\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__13070\,
            I => \N__13046\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13039\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13039\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13039\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13036\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13031\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13031\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__13049\,
            I => \N__13026\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__13046\,
            I => \N__13026\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13039\,
            I => \N__13023\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__13036\,
            I => \N__13020\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13031\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__13026\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__13023\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__13020\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__13011\,
            I => \N__13005\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13010\,
            I => \N__13002\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12995\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13008\,
            I => \N__12995\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12995\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13002\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__12995\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__12990\,
            I => \N__12987\
        );

    \I__2420\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12982\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12977\
        );

    \I__2418\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12977\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__12982\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__12977\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__2415\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12968\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__12971\,
            I => \N__12963\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__12968\,
            I => \N__12959\
        );

    \I__2412\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12956\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__12966\,
            I => \N__12953\
        );

    \I__2410\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12950\
        );

    \I__2409\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12947\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__12959\,
            I => \N__12944\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__12956\,
            I => \N__12941\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12938\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__12950\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__12947\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__12944\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__12941\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__12938\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__12927\,
            I => \N__12922\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12916\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12916\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12913\
        );

    \I__2396\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12908\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__12916\,
            I => \N__12905\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12913\,
            I => \N__12902\
        );

    \I__2393\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12897\
        );

    \I__2392\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12897\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12888\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__12905\,
            I => \N__12888\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__12902\,
            I => \N__12888\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12888\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__12888\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__2385\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12878\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__12881\,
            I => \N__12874\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__12878\,
            I => \N__12870\
        );

    \I__2382\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12865\
        );

    \I__2381\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12865\
        );

    \I__2380\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12862\
        );

    \I__2379\ : Span4Mux_s2_h
    port map (
            O => \N__12870\,
            I => \N__12857\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__12865\,
            I => \N__12857\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__12862\,
            I => \uu2.N_106\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__12857\,
            I => \uu2.N_106\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__12852\,
            I => \N__12846\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__12851\,
            I => \N__12843\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12839\
        );

    \I__2372\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12834\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12846\,
            I => \N__12834\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12843\,
            I => \N__12829\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12829\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__12839\,
            I => \N__12826\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__12834\,
            I => \N__12823\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__12829\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__12826\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__12823\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2363\ : CEMux
    port map (
            O => \N__12816\,
            I => \N__12812\
        );

    \I__2362\ : CEMux
    port map (
            O => \N__12815\,
            I => \N__12809\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__12812\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12809\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__12804\,
            I => \N__12801\
        );

    \I__2358\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__12798\,
            I => \G_193\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__12795\,
            I => \G_193_cascade_\
        );

    \I__2355\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12789\,
            I => \Lab_UT.dispString.N_219\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__12786\,
            I => \Lab_UT.dispString.N_222_cascade_\
        );

    \I__2352\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12780\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__12780\,
            I => \N__12776\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__12779\,
            I => \N__12773\
        );

    \I__2349\ : Span4Mux_s2_v
    port map (
            O => \N__12776\,
            I => \N__12770\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12767\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__12770\,
            I => \N__12761\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__12767\,
            I => \N__12761\
        );

    \I__2345\ : InMux
    port map (
            O => \N__12766\,
            I => \N__12758\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__12761\,
            I => \L3_tx_data_3\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__12758\,
            I => \L3_tx_data_3\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__12753\,
            I => \N__12750\
        );

    \I__2341\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12747\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__12747\,
            I => \G_189\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__12744\,
            I => \G_189_cascade_\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12738\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__12738\,
            I => \Lab_UT.dispString.un42_dOutP\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__2333\ : Span4Mux_s2_v
    port map (
            O => \N__12726\,
            I => \N__12722\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \N__12718\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__12722\,
            I => \N__12715\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12712\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12709\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__12715\,
            I => \L3_tx_data_6\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__12712\,
            I => \L3_tx_data_6\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12709\,
            I => \L3_tx_data_6\
        );

    \I__2325\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12698\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12695\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12698\,
            I => \N__12692\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__12695\,
            I => \N__12688\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__12692\,
            I => \N__12685\
        );

    \I__2320\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12682\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__12688\,
            I => \uu0_sec_clkD\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__12685\,
            I => \uu0_sec_clkD\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__12682\,
            I => \uu0_sec_clkD\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12672\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12672\,
            I => \Lab_UT.dispString.m44_ns_1\
        );

    \I__2314\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12657\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12657\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12657\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12657\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__12657\,
            I => \N__12654\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__12654\,
            I => \N__12648\
        );

    \I__2308\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12641\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12641\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12641\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__12648\,
            I => \Lab_UT.sec2_0\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12641\,
            I => \Lab_UT.sec2_0\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12632\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12629\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__12632\,
            I => \G_190\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__12629\,
            I => \G_190\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__12624\,
            I => \G_190_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12618\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__12618\,
            I => \Lab_UT.dispString.i21_mux\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__12615\,
            I => \Lab_UT.dispString.m28_ns_1_cascade_\
        );

    \I__2295\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12609\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12609\,
            I => \Lab_UT.dispString.N_204\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__12606\,
            I => \N__12601\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12596\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12596\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12593\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__12596\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12593\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2287\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12585\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__12585\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__12582\,
            I => \N__12575\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \N__12572\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12568\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__12579\,
            I => \N__12564\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12561\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12551\
        );

    \I__2279\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12551\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12551\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12548\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__12567\,
            I => \N__12544\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12541\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12561\,
            I => \N__12538\
        );

    \I__2273\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12531\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12531\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12531\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__12551\,
            I => \N__12528\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__12548\,
            I => \N__12525\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12520\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12520\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12541\,
            I => \N__12515\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__12538\,
            I => \N__12515\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12531\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__12528\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__12525\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12520\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__12515\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12501\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12501\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__12498\,
            I => \N__12495\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12492\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12492\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12483\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__12488\,
            I => \N__12480\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12476\
        );

    \I__2251\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12472\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__12483\,
            I => \N__12469\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12464\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12464\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12476\,
            I => \N__12461\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12458\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12472\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__12469\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12464\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__12461\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12458\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12444\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12444\,
            I => \uu2.bitmap_pmux_24_am_1\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12424\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12424\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12424\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12424\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12424\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12419\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12419\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12414\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__12419\,
            I => \N__12414\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__12414\,
            I => \Lab_UT.min1_1\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12408\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12408\,
            I => \N__12405\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__12405\,
            I => \Lab_UT.dispString.un46_dOutP_2\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12399\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12399\,
            I => \uu2.bitmap_pmux_24_bm_1\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12393\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__12393\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__12390\,
            I => \N__12387\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12384\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12384\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12378\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__12378\,
            I => \N__12370\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12363\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12363\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12363\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12355\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12352\
        );

    \I__2211\ : Span4Mux_v
    port map (
            O => \N__12370\,
            I => \N__12347\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12363\,
            I => \N__12347\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12344\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12341\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12338\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12333\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12333\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12355\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12352\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__12347\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12344\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__12341\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12338\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__12333\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2197\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12315\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__12312\,
            I => \N__12309\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__12309\,
            I => \uu2.bitmap_RNI5T9T1Z0Z_72\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12303\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__12300\,
            I => \uu2.bitmap_pmux_sn_N_54_mux\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12294\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12294\,
            I => \uu2.N_237\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12288\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12288\,
            I => \N__12285\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__12285\,
            I => \uu2.bitmap_pmux_sn_N_15\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__12282\,
            I => \uu2.N_395_cascade_\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12279\,
            I => \N__12276\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12276\,
            I => \N__12273\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__12273\,
            I => \uu2.N_401\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12267\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__12267\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12259\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__12263\,
            I => \N__12254\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12249\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12259\,
            I => \N__12246\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12243\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12234\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12234\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12234\
        );

    \I__2171\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12234\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12249\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12246\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__12243\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12234\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12219\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__12216\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12210\,
            I => \uu2.bitmap_pmux_15_i_m2_ns_1\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12204\,
            I => \uu2.N_123\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__12201\,
            I => \N__12196\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12187\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12184\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12180\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12177\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12168\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12168\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12168\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12168\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12165\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12160\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12160\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12157\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__12180\,
            I => \N__12154\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__12177\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12168\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12165\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__12160\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__12157\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__12154\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2138\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12138\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__12132\,
            I => \uu2.bitmap_RNIU2ISZ0Z_52\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12126\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12126\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2132\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__12120\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__12117\,
            I => \N__12114\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12111\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__12111\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12105\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12105\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12099\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12092\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12086\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12083\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12080\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12075\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12075\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12086\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__12083\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__12080\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12075\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12063\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__12060\,
            I => \N__12054\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12048\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12048\
        );

    \I__2108\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12045\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12040\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12040\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12048\,
            I => \N__12037\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__12045\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12040\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__12037\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__2101\ : CEMux
    port map (
            O => \N__12030\,
            I => \N__12027\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__12027\,
            I => \N__12022\
        );

    \I__2099\ : CEMux
    port map (
            O => \N__12026\,
            I => \N__12019\
        );

    \I__2098\ : CEMux
    port map (
            O => \N__12025\,
            I => \N__12016\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__12022\,
            I => \N__12011\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__12011\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__12016\,
            I => \N__12008\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__12011\,
            I => \N__12005\
        );

    \I__2093\ : Sp12to4
    port map (
            O => \N__12008\,
            I => \N__12002\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__12005\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__12002\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2090\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11994\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__11994\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__11991\,
            I => \N__11988\
        );

    \I__2087\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11983\
        );

    \I__2086\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11980\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11977\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11983\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__11980\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__11977\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2081\ : InMux
    port map (
            O => \N__11970\,
            I => \N__11966\
        );

    \I__2080\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11963\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__11966\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__11963\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11954\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__11957\,
            I => \N__11951\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11948\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11945\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__11948\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11945\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2071\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11935\
        );

    \I__2070\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11930\
        );

    \I__2069\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11930\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__11935\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__11930\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__2065\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11915\
        );

    \I__2064\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11915\
        );

    \I__2063\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11912\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__11915\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__11912\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__11907\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__11904\,
            I => \N__11901\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11892\
        );

    \I__2056\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11887\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11887\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__11895\,
            I => \N__11884\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__11892\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__11887\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__11884\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11874\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__11874\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__11871\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11861\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11858\
        );

    \I__2045\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11851\
        );

    \I__2044\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11851\
        );

    \I__2043\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11851\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__11861\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__11858\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__11851\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2039\ : IoInMux
    port map (
            O => \N__11844\,
            I => \N__11841\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__11841\,
            I => \N__11838\
        );

    \I__2037\ : IoSpan4Mux
    port map (
            O => \N__11838\,
            I => \N__11835\
        );

    \I__2036\ : Span4Mux_s1_v
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__11832\,
            I => \buart.Z_rx.sample\
        );

    \I__2034\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11814\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11814\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11811\
        );

    \I__2031\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11804\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11804\
        );

    \I__2029\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11804\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11797\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11797\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11797\
        );

    \I__2025\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11791\
        );

    \I__2024\ : InMux
    port map (
            O => \N__11819\,
            I => \N__11791\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__11814\,
            I => \N__11782\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__11811\,
            I => \N__11782\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11804\,
            I => \N__11782\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__11797\,
            I => \N__11782\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11779\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11791\,
            I => \buart.Z_rx.startbit\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__11782\,
            I => \buart.Z_rx.startbit\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__11779\,
            I => \buart.Z_rx.startbit\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__11772\,
            I => \N__11768\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__11771\,
            I => \N__11765\
        );

    \I__2013\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11760\
        );

    \I__2012\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11753\
        );

    \I__2011\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11753\
        );

    \I__2010\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11753\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__11760\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__11753\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \buart.Z_rx.idle_0_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11740\
        );

    \I__2005\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11737\
        );

    \I__2004\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11734\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__11740\,
            I => \N__11731\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__11737\,
            I => \buart.Z_rx.idle\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__11734\,
            I => \buart.Z_rx.idle\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__11731\,
            I => \buart.Z_rx.idle\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__1998\ : InMux
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__11715\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \N__11708\
        );

    \I__1994\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11702\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11699\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11692\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11692\
        );

    \I__1990\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11692\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__11702\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__11699\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11692\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__11685\,
            I => \N__11682\
        );

    \I__1985\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11675\
        );

    \I__1984\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11672\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11669\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11664\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11664\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__11675\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__11672\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__11669\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__11664\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__11655\,
            I => \N__11652\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11646\
        );

    \I__1974\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11643\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11638\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11638\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__11646\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__11643\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__11638\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__11631\,
            I => \buart.Z_rx.valid_1_cascade_\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11621\
        );

    \I__1966\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11618\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11611\
        );

    \I__1964\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11611\
        );

    \I__1963\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11611\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__11621\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11618\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__11611\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__11604\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11597\
        );

    \I__1957\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11594\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11589\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__11594\,
            I => \N__11589\
        );

    \I__1954\ : Odrv12
    port map (
            O => \N__11589\,
            I => \Lab_UT.dispString.N_191\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__11583\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2\
        );

    \I__1951\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11576\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11573\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__11576\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__11573\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11568\,
            I => \N__11565\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11565\,
            I => \buart.Z_tx.uart_busy_0_0\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11559\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__11559\,
            I => \N__11555\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11552\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__11555\,
            I => \N__11549\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11552\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__11549\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1939\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11533\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11533\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11533\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11528\
        );

    \I__1935\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11528\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__11533\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11528\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \N__11520\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11511\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11511\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11504\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11504\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11504\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11511\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11504\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11495\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__11498\,
            I => \N__11491\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11484\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11484\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11484\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__11484\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__11481\,
            I => \N__11476\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11472\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11467\
        );

    \I__1915\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11467\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11464\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__11472\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11467\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__11464\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1910\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__11454\,
            I => \buart.Z_tx.un1_bitcount_c3\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11448\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11448\,
            I => vbuf_tx_data_0
        );

    \I__1906\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11442\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11436\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1902\ : IoInMux
    port map (
            O => \N__11433\,
            I => \N__11430\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11430\,
            I => \N__11427\
        );

    \I__1900\ : Span4Mux_s3_h
    port map (
            O => \N__11427\,
            I => \N__11424\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__11424\,
            I => \N__11421\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__11421\,
            I => o_serial_data_c
        );

    \I__1897\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11415\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11415\,
            I => vbuf_tx_data_1
        );

    \I__1895\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11409\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11409\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11403\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11403\,
            I => vbuf_tx_data_2
        );

    \I__1891\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11397\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11397\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11391\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__11391\,
            I => vbuf_tx_data_3
        );

    \I__1887\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11385\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1885\ : InMux
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__11379\,
            I => vbuf_tx_data_4
        );

    \I__1883\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11373\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__11373\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11367\,
            I => vbuf_tx_data_5
        );

    \I__1879\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11361\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \Lab_UT.dispString.N_211_cascade_\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11352\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_2\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11346\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__11346\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_2\
        );

    \I__1872\ : CEMux
    port map (
            O => \N__11343\,
            I => \N__11340\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11340\,
            I => \N__11337\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__11337\,
            I => \N__11334\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__11334\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11325\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__11322\,
            I => \N__11317\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11314\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11311\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__11317\,
            I => \L3_tx_data_4\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11314\,
            I => \L3_tx_data_4\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11311\,
            I => \L3_tx_data_4\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11304\,
            I => \N__11299\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11296\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11293\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__11299\,
            I => \L3_tx_data_2\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11296\,
            I => \L3_tx_data_2\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11293\,
            I => \L3_tx_data_2\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__11286\,
            I => \uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11280\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11280\,
            I => \N__11277\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__11277\,
            I => \N__11272\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11269\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11266\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__11272\,
            I => \L3_tx_data_0\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11269\,
            I => \L3_tx_data_0\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11266\,
            I => \L3_tx_data_0\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11241\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11241\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11241\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11241\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11236\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11236\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11253\,
            I => \N__11233\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11230\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11225\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11225\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11241\,
            I => \N__11220\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11220\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11217\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11214\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11225\,
            I => \N__11211\
        );

    \I__1829\ : Span4Mux_s2_h
    port map (
            O => \N__11220\,
            I => \N__11208\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11217\,
            I => \N__11200\
        );

    \I__1827\ : Span4Mux_h
    port map (
            O => \N__11214\,
            I => \N__11197\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__11211\,
            I => \N__11194\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__11208\,
            I => \N__11191\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11186\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11186\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11179\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11179\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11179\
        );

    \I__1819\ : Odrv12
    port map (
            O => \N__11200\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__11197\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__11194\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__11191\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11186\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__11179\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__11166\,
            I => \N__11163\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11160\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11157\
        );

    \I__1810\ : Span12Mux_s6_v
    port map (
            O => \N__11157\,
            I => \N__11152\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11149\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11146\
        );

    \I__1807\ : Odrv12
    port map (
            O => \N__11152\,
            I => \L3_tx_data_5\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11149\,
            I => \L3_tx_data_5\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11146\,
            I => \L3_tx_data_5\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__11139\,
            I => \Lab_UT.didp.countrce1.q_5_0_cascade_\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11133\,
            I => \N__11121\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11121\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11121\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11121\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11121\,
            I => \N__11115\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11108\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11108\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11118\,
            I => \N__11108\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__11115\,
            I => \Lab_UT.sec2_1\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11108\,
            I => \Lab_UT.sec2_1\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11091\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11091\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11091\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11091\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11091\,
            I => \N__11086\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__11090\,
            I => \N__11083\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11089\,
            I => \N__11080\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__11086\,
            I => \N__11076\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11069\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11069\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11069\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__11076\,
            I => \Lab_UT.sec2_2\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11069\,
            I => \Lab_UT.sec2_2\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__11064\,
            I => \N__11057\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11054\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__11062\,
            I => \N__11051\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11046\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11037\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11037\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11037\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11037\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11030\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11030\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11030\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__11027\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__11027\,
            I => \Lab_UT.sec2_3\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__11024\,
            I => \Lab_UT.sec2_3\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__11013\,
            I => \uu2.un28_w_addr_user_i_0_a2_0Z0Z_4\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__11010\,
            I => \Lab_UT.dispString.un42_dOutP_cascade_\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__11004\,
            I => \uu2.un28_w_addr_user_i_0_a2_0Z0Z_0\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__1757\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__10995\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__1755\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__10989\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__1753\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__10983\,
            I => \uu2.bitmap_pmux_25_i_m2_bm_1\
        );

    \I__1751\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10974\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10971\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10965\
        );

    \I__1748\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10965\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10960\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10960\
        );

    \I__1745\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10957\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__10965\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__10960\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10957\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__10950\,
            I => \uu2.bitmap_pmux_21_ns_1_cascade_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10944\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__10944\,
            I => \N__10941\
        );

    \I__1738\ : Span4Mux_h
    port map (
            O => \N__10941\,
            I => \N__10938\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__10938\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__10935\,
            I => \uu2.N_393_cascade_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__10929\,
            I => \uu2.N_397\
        );

    \I__1733\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10920\
        );

    \I__1732\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10920\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__10920\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__1730\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10914\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__10914\,
            I => \uu2.N_128\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10908\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__10908\,
            I => \uu2.N_131\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10902\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10899\
        );

    \I__1724\ : Span4Mux_h
    port map (
            O => \N__10899\,
            I => \N__10895\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10892\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__10895\,
            I => \N__10887\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__10892\,
            I => \N__10887\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__10887\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__10881\,
            I => \uu2.bitmap_RNIFJI02Z0Z_212\
        );

    \I__1717\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10871\
        );

    \I__1716\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10871\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10868\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10865\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__10868\,
            I => \N__10862\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__10865\,
            I => \uu2.N_65\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__10862\,
            I => \uu2.N_65\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10854\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__10854\,
            I => \N__10851\
        );

    \I__1708\ : Odrv12
    port map (
            O => \N__10851\,
            I => \uu2.bitmap_pmux_u_0_83_0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10832\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10832\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10832\
        );

    \I__1704\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10832\
        );

    \I__1703\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10832\
        );

    \I__1702\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10824\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__10832\,
            I => \N__10821\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10818\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10809\
        );

    \I__1698\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10809\
        );

    \I__1697\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10809\
        );

    \I__1696\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10809\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10824\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__10821\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__10818\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__10809\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__10799\,
            I => \N__10790\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__10798\,
            I => \N__10784\
        );

    \I__1688\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10780\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10771\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10771\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10771\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10789\,
            I => \N__10771\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10764\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10764\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10784\,
            I => \N__10764\
        );

    \I__1680\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10761\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__10780\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__10771\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__10764\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__10761\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__1675\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10749\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10749\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10743\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10743\,
            I => \uu2.N_112_i\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__10740\,
            I => \uu2.N_100_cascade_\
        );

    \I__1670\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10734\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10734\,
            I => \uu2.N_921_tz_tz\
        );

    \I__1668\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__10728\,
            I => \N__10725\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__10725\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__10722\,
            I => \uu2.N_923_tz_cascade_\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__10713\,
            I => \uu2.w_addr_displaying_RNI8ND5GZ0Z_3\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__10710\,
            I => \N__10707\
        );

    \I__1660\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1659\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10701\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10692\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10687\
        );

    \I__1656\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10687\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10675\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10675\
        );

    \I__1653\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10675\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10675\
        );

    \I__1651\ : Span12Mux_s4_h
    port map (
            O => \N__10692\,
            I => \N__10672\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10687\,
            I => \N__10669\
        );

    \I__1649\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10662\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10662\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10662\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__10675\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__10672\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1644\ : Odrv12
    port map (
            O => \N__10669\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__10662\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__10653\,
            I => \N__10650\
        );

    \I__1641\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10645\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__10649\,
            I => \N__10642\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__10648\,
            I => \N__10639\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__10645\,
            I => \N__10633\
        );

    \I__1637\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10624\
        );

    \I__1636\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10624\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10624\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10624\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10621\
        );

    \I__1632\ : Span4Mux_s1_v
    port map (
            O => \N__10633\,
            I => \N__10618\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__10624\,
            I => \N__10615\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__10621\,
            I => \N__10612\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__10618\,
            I => \uu2.N_34\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__10615\,
            I => \uu2.N_34\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__10612\,
            I => \uu2.N_34\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10601\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \N__10597\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__10601\,
            I => \N__10592\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10587\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10587\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__10596\,
            I => \N__10583\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10580\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__10592\,
            I => \N__10574\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10587\,
            I => \N__10574\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10569\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10566\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__10580\,
            I => \N__10563\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10560\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__10574\,
            I => \N__10557\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10552\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10552\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__10569\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__10566\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__10563\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10560\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__10557\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10552\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__10536\,
            I => \N__10533\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__10533\,
            I => \N__10530\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__10530\,
            I => \uu2.N_47\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__10526\,
            I => \N__10518\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__10525\,
            I => \N__10514\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10502\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10502\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10502\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10502\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10502\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10499\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10496\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10499\,
            I => \N__10493\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__10496\,
            I => \N__10490\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__10493\,
            I => \uu2.N_38\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__10490\,
            I => \uu2.N_38\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10473\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10456\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10456\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10456\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10456\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10456\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10456\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10456\
        );

    \I__1578\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10456\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10453\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10448\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10448\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10445\
        );

    \I__1573\ : Span4Mux_s1_v
    port map (
            O => \N__10448\,
            I => \N__10442\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__10445\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_5\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__10442\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_5\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10428\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10428\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10428\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10417\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10417\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10414\
        );

    \I__1563\ : Span4Mux_s3_h
    port map (
            O => \N__10422\,
            I => \N__10409\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10409\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10414\,
            I => \uu2.N_33\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__10409\,
            I => \uu2.N_33\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10392\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10392\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10392\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10384\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10384\
        );

    \I__1554\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10384\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10392\,
            I => \N__10381\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10371\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10384\,
            I => \N__10368\
        );

    \I__1550\ : Span4Mux_h
    port map (
            O => \N__10381\,
            I => \N__10365\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10362\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10357\
        );

    \I__1547\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10357\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10348\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10348\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10348\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10348\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10371\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__10368\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__10365\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10362\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10357\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10348\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10325\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10321\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__10333\,
            I => \N__10318\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10313\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10310\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10303\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10303\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10303\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10298\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10298\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10294\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10291\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10286\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10286\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10283\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10276\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10276\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__10298\,
            I => \N__10276\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10270\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10294\,
            I => \N__10265\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10291\,
            I => \N__10265\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10258\
        );

    \I__1514\ : Span4Mux_h
    port map (
            O => \N__10283\,
            I => \N__10258\
        );

    \I__1513\ : Span4Mux_s3_h
    port map (
            O => \N__10276\,
            I => \N__10258\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10255\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10250\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10250\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10270\,
            I => \L3_tx_data_rdy\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__10265\,
            I => \L3_tx_data_rdy\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__10258\,
            I => \L3_tx_data_rdy\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__10255\,
            I => \L3_tx_data_rdy\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10250\,
            I => \L3_tx_data_rdy\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__10230\,
            I => \uu2.mem0.N_136\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10224\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10224\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10218\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__10215\,
            I => \uu2.bitmap_pmux_25_i_m2_am_1_cascade_\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__10206\,
            I => \uu2.bitmap_RNIG91I1Z0Z_66\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10197\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10197\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__1489\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10191\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10191\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10185\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__10185\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10179\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10176\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10170\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10170\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10167\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10164\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10161\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10158\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10155\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10152\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10149\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__10140\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10133\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10130\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10130\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__10127\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__10122\,
            I => \N__10118\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10111\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10108\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10103\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10103\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10098\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10098\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10111\,
            I => \N__10095\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10092\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10103\,
            I => \N__10089\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10086\
        );

    \I__1454\ : Span4Mux_s3_h
    port map (
            O => \N__10095\,
            I => \N__10083\
        );

    \I__1453\ : Span4Mux_s2_h
    port map (
            O => \N__10092\,
            I => \N__10080\
        );

    \I__1452\ : Span12Mux_s3_h
    port map (
            O => \N__10089\,
            I => \N__10077\
        );

    \I__1451\ : Span4Mux_s3_h
    port map (
            O => \N__10086\,
            I => \N__10074\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__10083\,
            I => \N__10071\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__10080\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__10077\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__10074\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__10071\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10058\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10055\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10058\,
            I => \N__10052\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10055\,
            I => \N__10046\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__10052\,
            I => \N__10043\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10036\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10036\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10036\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__10046\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__10043\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10036\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10024\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10021\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10018\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10015\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10021\,
            I => \N__10012\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10018\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__10015\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__10012\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9998\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9998\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10003\,
            I => \N__9995\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9992\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__9995\,
            I => \N__9989\
        );

    \I__1421\ : Span4Mux_s3_h
    port map (
            O => \N__9992\,
            I => \N__9986\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__9989\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__9986\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9978\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__9978\,
            I => \N__9975\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__9972\,
            I => \uu2.mem0.N_54_i\
        );

    \I__1414\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9966\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9963\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__9963\,
            I => \N__9960\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__9960\,
            I => \uu2.r_data_wire_0\
        );

    \I__1410\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__9954\,
            I => \N__9951\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__9948\,
            I => \uu2.r_data_wire_1\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9942\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__9939\,
            I => \N__9936\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__9936\,
            I => \uu2.r_data_wire_2\
        );

    \I__1402\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9930\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__9930\,
            I => \N__9927\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__9927\,
            I => \N__9924\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__9924\,
            I => \uu2.r_data_wire_3\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9918\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__9918\,
            I => \N__9915\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__9915\,
            I => \N__9912\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__9912\,
            I => \uu2.r_data_wire_4\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9906\,
            I => \N__9903\
        );

    \I__1392\ : Span4Mux_v
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__9900\,
            I => \uu2.r_data_wire_5\
        );

    \I__1390\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__9891\,
            I => \N__9888\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__9888\,
            I => \uu2.r_data_wire_6\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__9882\,
            I => \N__9879\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9876\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__9876\,
            I => \uu2.r_data_wire_7\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__9873\,
            I => \uu2.N_106_cascade_\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__9870\,
            I => \N__9867\
        );

    \I__1380\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9861\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__9861\,
            I => \uu2.N_164\
        );

    \I__1377\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9854\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__9857\,
            I => \N__9851\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9847\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9840\
        );

    \I__1373\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9840\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__9847\,
            I => \N__9837\
        );

    \I__1371\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9832\
        );

    \I__1370\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9832\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__9840\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__9837\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__9832\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9822\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9822\,
            I => \uu2.w_addr_user_3_i_a2_3_6\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__9819\,
            I => \uu2.w_addr_user_3_i_a2_2_6_cascade_\
        );

    \I__1363\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9811\
        );

    \I__1362\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9808\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9805\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9811\,
            I => \uu2.N_230\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__9808\,
            I => \uu2.N_230\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__9805\,
            I => \uu2.N_230\
        );

    \I__1357\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9792\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9789\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9784\
        );

    \I__1354\ : InMux
    port map (
            O => \N__9795\,
            I => \N__9784\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__9792\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__9789\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__9784\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__1347\ : Span4Mux_s3_h
    port map (
            O => \N__9768\,
            I => \N__9765\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__9765\,
            I => \uu2.mem0.N_138\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__9762\,
            I => \oneSecStrb_cascade_\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__9759\,
            I => \N__9755\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9752\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__9755\,
            I => \N__9749\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9746\
        );

    \I__1340\ : Span12Mux_s9_v
    port map (
            O => \N__9749\,
            I => \N__9741\
        );

    \I__1339\ : Span12Mux_s5_h
    port map (
            O => \N__9746\,
            I => \N__9741\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__9741\,
            I => clk
        );

    \I__1337\ : SRMux
    port map (
            O => \N__9738\,
            I => \N__9734\
        );

    \I__1336\ : CEMux
    port map (
            O => \N__9737\,
            I => \N__9731\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9728\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9731\,
            I => \N__9725\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__9728\,
            I => \N__9720\
        );

    \I__1332\ : Span4Mux_h
    port map (
            O => \N__9725\,
            I => \N__9720\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__9720\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__9717\,
            I => \N__9711\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9706\
        );

    \I__1328\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9701\
        );

    \I__1327\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9701\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9694\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9694\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9694\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9691\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9686\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__9694\,
            I => \N__9686\
        );

    \I__1320\ : Span4Mux_s3_h
    port map (
            O => \N__9691\,
            I => \N__9682\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__9686\,
            I => \N__9679\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9676\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__9682\,
            I => \N__9673\
        );

    \I__1316\ : Span4Mux_s2_v
    port map (
            O => \N__9679\,
            I => \N__9668\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__9676\,
            I => \N__9668\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__9673\,
            I => \uu2.N_102\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__9668\,
            I => \uu2.N_102\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__9663\,
            I => \N__9658\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9655\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9650\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9650\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__9655\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__9650\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__9645\,
            I => \uu2.N_161_cascade_\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__9642\,
            I => \uu2.N_101_cascade_\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__9639\,
            I => \N__9633\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \N__9628\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__9637\,
            I => \N__9625\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9618\
        );

    \I__1300\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9618\
        );

    \I__1299\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9618\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__9631\,
            I => \N__9615\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9612\
        );

    \I__1296\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9609\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9606\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9603\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__9612\,
            I => \N__9600\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9609\,
            I => \N__9597\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__9606\,
            I => \N__9594\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__9603\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1289\ : Odrv12
    port map (
            O => \N__9600\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__9597\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__9594\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__9585\,
            I => \N__9581\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9578\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9575\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9571\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9568\
        );

    \I__1281\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9561\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__9571\,
            I => \N__9556\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__9568\,
            I => \N__9556\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9547\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9547\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9547\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9547\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__9561\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__9556\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9547\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__9540\,
            I => \N__9537\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__9531\,
            I => \uu2.mem0.N_135\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__9522\,
            I => \uu2.mem0.N_134\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__9519\,
            I => \uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_\
        );

    \I__1263\ : CEMux
    port map (
            O => \N__9516\,
            I => \N__9512\
        );

    \I__1262\ : CEMux
    port map (
            O => \N__9515\,
            I => \N__9509\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9506\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9509\,
            I => \N__9503\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__9506\,
            I => \N__9500\
        );

    \I__1258\ : Span4Mux_s0_v
    port map (
            O => \N__9503\,
            I => \N__9497\
        );

    \I__1257\ : Span4Mux_s0_h
    port map (
            O => \N__9500\,
            I => \N__9494\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__9497\,
            I => \uu2.N_32_0\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__9494\,
            I => \uu2.N_32_0\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__9480\,
            I => \uu2.mem0.N_133\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__9477\,
            I => \N__9471\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9459\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9459\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9459\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9459\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9459\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9459\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9453\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9453\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9447\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9441\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__1236\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9432\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__9429\,
            I => \uu2.bitmap_RNIRETJ1Z0Z_93_cascade_\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__9426\,
            I => \uu2.bitmap_pmux_27_ns_1_cascade_\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9417\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9414\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__9414\,
            I => \uu2.N_404\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9408\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__1226\ : Span4Mux_s3_h
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__9402\,
            I => \uu2.bitmap_pmux_u_0_a2_0_2_0\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9394\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9389\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9389\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N__9385\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9382\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__9388\,
            I => \N__9377\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__9385\,
            I => \N__9371\
        );

    \I__1217\ : Span4Mux_s3_h
    port map (
            O => \N__9382\,
            I => \N__9368\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9359\
        );

    \I__1215\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9359\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9359\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9359\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9354\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9354\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__9371\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__9368\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__9359\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9354\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__9345\,
            I => \uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9335\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9328\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9328\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9328\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9325\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9335\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9328\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9325\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9304\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9304\
        );

    \I__1195\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9304\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9304\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9299\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9299\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9304\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9299\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__9294\,
            I => \N__9290\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__9293\,
            I => \N__9287\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9283\
        );

    \I__1186\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9280\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9277\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9283\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9280\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__9277\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__9270\,
            I => \N__9264\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9259\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9259\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9256\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9253\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9250\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__9256\,
            I => \uu2.un306_ci\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9253\,
            I => \uu2.un306_ci\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__9250\,
            I => \uu2.un306_ci\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9236\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9236\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9233\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9236\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9233\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__9228\,
            I => \uu2.un306_ci_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9216\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9216\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9211\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9211\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9208\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9216\,
            I => \N__9203\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__9211\,
            I => \N__9203\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9208\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__9203\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9194\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9191\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9194\,
            I => \uu2.un284_ci\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9191\,
            I => \uu2.un284_ci\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__9186\,
            I => \N__9181\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9172\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9172\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9172\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9169\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9166\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9163\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9169\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9166\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__9163\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9152\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9149\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9152\,
            I => \uu2.un350_ci\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9149\,
            I => \uu2.un350_ci\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__9144\,
            I => \N__9140\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9134\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9134\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9131\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__9134\,
            I => \N__9128\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9131\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__9128\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9119\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9116\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9113\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9110\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9106\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9103\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9100\
        );

    \I__1125\ : Span4Mux_v
    port map (
            O => \N__9106\,
            I => \N__9095\
        );

    \I__1124\ : Span4Mux_h
    port map (
            O => \N__9103\,
            I => \N__9095\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9100\,
            I => \uu0.un88_ci_3\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__9095\,
            I => \uu0.un88_ci_3\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9081\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9078\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9075\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9072\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__9081\,
            I => \N__9067\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9067\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9075\,
            I => \N__9064\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9072\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__9067\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__9064\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9051\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__9048\
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__9048\,
            I => \uu0.un99_ci_0\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__9045\,
            I => \uu2.w_data_0_a2_0_6_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9034\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9023\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9023\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9023\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9023\
        );

    \I__1100\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9023\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9034\,
            I => \N__9018\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__9023\,
            I => \N__9018\
        );

    \I__1097\ : Span4Mux_v
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__9015\,
            I => \uu2.w_data_0_a2_2_6\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__9012\,
            I => \uu2.un1_l_count_2_2_cascade_\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__9009\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9006\,
            I => \N__9000\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9000\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9000\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8992\
        );

    \I__1089\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8987\
        );

    \I__1088\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8987\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__8992\,
            I => \N__8984\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__8987\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__8984\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__8979\,
            I => \N__8974\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \N__8971\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__8977\,
            I => \N__8968\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8961\
        );

    \I__1080\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8961\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8961\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__8961\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__1077\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__8955\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__1075\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8946\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8943\
        );

    \I__1073\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8940\
        );

    \I__1072\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8937\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8933\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__8943\,
            I => \N__8930\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__8940\,
            I => \N__8927\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__8937\,
            I => \N__8924\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8921\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__8933\,
            I => \uu0.un66_ci\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__8930\,
            I => \uu0.un66_ci\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__8927\,
            I => \uu0.un66_ci\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__8924\,
            I => \uu0.un66_ci\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__8921\,
            I => \uu0.un66_ci\
        );

    \I__1061\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8905\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8900\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8900\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8893\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8893\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__8899\,
            I => \N__8890\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__8898\,
            I => \N__8886\
        );

    \I__1054\ : Span4Mux_v
    port map (
            O => \N__8893\,
            I => \N__8879\
        );

    \I__1053\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8876\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8871\
        );

    \I__1051\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8871\
        );

    \I__1050\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8862\
        );

    \I__1049\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8862\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8862\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8862\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__8879\,
            I => \uu0.un110_ci\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__8876\,
            I => \uu0.un110_ci\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8871\,
            I => \uu0.un110_ci\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8862\,
            I => \uu0.un110_ci\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8844\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8844\
        );

    \I__1040\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8844\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__8841\,
            I => \uu0.un198_ci_2\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__8838\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8825\
        );

    \I__1035\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8825\
        );

    \I__1034\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8825\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8822\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8825\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__8822\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8810\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8806\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8797\
        );

    \I__1027\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8790\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8790\
        );

    \I__1025\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8790\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8787\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8784\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8777\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8777\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8777\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8774\
        );

    \I__1018\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8771\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8768\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8763\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8763\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__8787\,
            I => \N__8758\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__8784\,
            I => \N__8758\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__8777\,
            I => \uu0.un4_l_count_0\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__8774\,
            I => \uu0.un4_l_count_0\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__8771\,
            I => \uu0.un4_l_count_0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__8768\,
            I => \uu0.un4_l_count_0\
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__8763\,
            I => \uu0.un4_l_count_0\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__8758\,
            I => \uu0.un4_l_count_0\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__8745\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8738\
        );

    \I__1004\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8735\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__8738\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__8735\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1001\ : CEMux
    port map (
            O => \N__8730\,
            I => \N__8709\
        );

    \I__1000\ : CEMux
    port map (
            O => \N__8729\,
            I => \N__8709\
        );

    \I__999\ : CEMux
    port map (
            O => \N__8728\,
            I => \N__8709\
        );

    \I__998\ : CEMux
    port map (
            O => \N__8727\,
            I => \N__8709\
        );

    \I__997\ : CEMux
    port map (
            O => \N__8726\,
            I => \N__8709\
        );

    \I__996\ : CEMux
    port map (
            O => \N__8725\,
            I => \N__8709\
        );

    \I__995\ : CEMux
    port map (
            O => \N__8724\,
            I => \N__8709\
        );

    \I__994\ : GlobalMux
    port map (
            O => \N__8709\,
            I => \N__8706\
        );

    \I__993\ : gio2CtrlBuf
    port map (
            O => \N__8706\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__8703\,
            I => \N__8697\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__8702\,
            I => \N__8694\
        );

    \I__990\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8684\
        );

    \I__989\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8684\
        );

    \I__988\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8684\
        );

    \I__987\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8684\
        );

    \I__986\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8681\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__8684\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__8681\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__983\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8669\
        );

    \I__982\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8669\
        );

    \I__981\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8666\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__8666\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__8663\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__8658\,
            I => \N__8654\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__8657\,
            I => \N__8650\
        );

    \I__975\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8643\
        );

    \I__974\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8643\
        );

    \I__973\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8643\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__8643\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__971\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8633\
        );

    \I__970\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8633\
        );

    \I__969\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8630\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8633\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8630\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__966\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__8622\,
            I => \uu0.un4_l_count_12\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__963\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8608\
        );

    \I__961\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8600\
        );

    \I__960\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8600\
        );

    \I__959\ : Span4Mux_h
    port map (
            O => \N__8608\,
            I => \N__8597\
        );

    \I__958\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8594\
        );

    \I__957\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8589\
        );

    \I__956\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8589\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__8600\,
            I => \N__8586\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__8597\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__8594\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__8589\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__8586\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__949\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8566\
        );

    \I__947\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8559\
        );

    \I__946\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8559\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__8566\,
            I => \N__8556\
        );

    \I__944\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8553\
        );

    \I__943\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8550\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8547\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__8556\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8553\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8550\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__8547\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__936\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8529\
        );

    \I__935\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8526\
        );

    \I__934\ : InMux
    port map (
            O => \N__8533\,
            I => \N__8520\
        );

    \I__933\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8520\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8517\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8514\
        );

    \I__930\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8511\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8508\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__8517\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__8514\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__8511\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__8508\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__924\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8493\
        );

    \I__923\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8490\
        );

    \I__922\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8485\
        );

    \I__921\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8485\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8480\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8480\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8485\,
            I => \uu2.un404_ci\
        );

    \I__917\ : Odrv12
    port map (
            O => \N__8480\,
            I => \uu2.un404_ci\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__915\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8468\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__8471\,
            I => \N__8465\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8461\
        );

    \I__912\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8455\
        );

    \I__911\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8455\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__8461\,
            I => \N__8452\
        );

    \I__909\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8449\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8446\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__8452\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__8449\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__905\ : Odrv12
    port map (
            O => \N__8446\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__8439\,
            I => \uu2.un404_ci_cascade_\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__902\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8429\
        );

    \I__901\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8429\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8426\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__898\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8418\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8418\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__8415\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__894\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8404\
        );

    \I__893\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8401\
        );

    \I__892\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8398\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__8404\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8401\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__8398\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__888\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8388\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8388\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__885\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8376\
        );

    \I__884\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8373\
        );

    \I__883\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8368\
        );

    \I__882\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8368\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8376\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8373\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8368\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__877\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8353\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__8357\,
            I => \N__8350\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__8356\,
            I => \N__8347\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8353\,
            I => \N__8344\
        );

    \I__873\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8339\
        );

    \I__872\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8339\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__8344\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8339\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__869\ : CEMux
    port map (
            O => \N__8334\,
            I => \N__8331\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__8331\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__866\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8319\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__8324\,
            I => \N__8316\
        );

    \I__864\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8311\
        );

    \I__863\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8311\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8319\,
            I => \N__8308\
        );

    \I__861\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8305\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8302\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__8308\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8305\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__8302\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__856\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8292\,
            I => \uu2.mem0.N_31_i\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__8289\,
            I => \uu2.mem0.N_61_cascade_\
        );

    \I__853\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8283\,
            I => \uu2.mem0.w_data_1\
        );

    \I__851\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8277\,
            I => \uu2.mem0.w_data_4\
        );

    \I__849\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8271\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8271\,
            I => \uu2.N_922_tz_tz\
        );

    \I__847\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8265\,
            I => \uu2.bitmap_pmux\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__8262\,
            I => \uu2.bitmap_pmux_cascade_\
        );

    \I__844\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8256\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__8256\,
            I => \uu2.mem0.w_data_3\
        );

    \I__842\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8249\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__8252\,
            I => \N__8246\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8243\
        );

    \I__839\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8240\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__8243\,
            I => \uu2.N_37\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8240\,
            I => \uu2.N_37\
        );

    \I__836\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8232\,
            I => \uu2.mem0.N_59\
        );

    \I__834\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__8226\,
            I => \uu2.mem0.w_data_0\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__8223\,
            I => \N__8218\
        );

    \I__831\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8208\
        );

    \I__830\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8208\
        );

    \I__829\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8208\
        );

    \I__828\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8208\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8208\,
            I => \uu0.un154_ci_9\
        );

    \I__826\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8200\
        );

    \I__825\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8195\
        );

    \I__824\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8195\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8200\,
            I => \N__8192\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8195\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__8192\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__8187\,
            I => \uu0.un4_l_count_0_8_cascade_\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__8184\,
            I => \N__8178\
        );

    \I__818\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8175\
        );

    \I__817\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8170\
        );

    \I__816\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8170\
        );

    \I__815\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8167\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8175\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8170\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8167\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__811\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8154\
        );

    \I__810\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8151\
        );

    \I__809\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8148\
        );

    \I__808\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8145\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8154\,
            I => \N__8140\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8151\,
            I => \N__8140\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8148\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8145\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__8140\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__802\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8128\
        );

    \I__801\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8125\
        );

    \I__800\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8122\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8128\,
            I => \N__8119\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8125\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8122\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__8119\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__8112\,
            I => \uu2.N_34_cascade_\
        );

    \I__794\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8106\,
            I => \uu2.N_114\
        );

    \I__792\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__8097\,
            I => \uu2.mem0.w_data_6\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__788\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8085\
        );

    \I__787\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8078\
        );

    \I__786\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8078\
        );

    \I__785\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8078\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8085\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8078\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__782\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__8067\,
            I => \uu0.un143_ci_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8046\
        );

    \I__778\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8046\
        );

    \I__777\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8046\
        );

    \I__776\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8046\
        );

    \I__775\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8046\
        );

    \I__774\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8046\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8046\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__8043\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__8040\,
            I => \N__8037\
        );

    \I__770\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8034\,
            I => \uu0.un165_ci_0\
        );

    \I__768\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8025\
        );

    \I__767\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8025\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8025\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__765\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8013\
        );

    \I__764\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8013\
        );

    \I__763\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8013\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8013\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__761\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8005\
        );

    \I__760\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8000\
        );

    \I__759\ : InMux
    port map (
            O => \N__8008\,
            I => \N__8000\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8005\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8000\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__7995\,
            I => \uu0.un55_ci_cascade_\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__7992\,
            I => \N__7985\
        );

    \I__754\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7971\
        );

    \I__753\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7971\
        );

    \I__752\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7971\
        );

    \I__751\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7971\
        );

    \I__750\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7971\
        );

    \I__749\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7971\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__7971\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__747\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7955\
        );

    \I__746\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7955\
        );

    \I__745\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7955\
        );

    \I__744\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7955\
        );

    \I__743\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7952\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__7955\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__7952\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__7947\,
            I => \N__7943\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__7946\,
            I => \N__7940\
        );

    \I__738\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7931\
        );

    \I__737\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7931\
        );

    \I__736\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7931\
        );

    \I__735\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7928\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__7931\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__7928\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7918\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7912\
        );

    \I__730\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7909\
        );

    \I__729\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7906\
        );

    \I__728\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7897\
        );

    \I__727\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7897\
        );

    \I__726\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7897\
        );

    \I__725\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7897\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__7909\,
            I => \N__7894\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7906\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__7897\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__7894\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__7887\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__719\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__7878\,
            I => \uu0.un4_l_count_18\
        );

    \I__716\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7870\
        );

    \I__715\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7865\
        );

    \I__714\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7865\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__7870\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__7865\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__7860\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__710\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7846\
        );

    \I__709\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7846\
        );

    \I__708\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7846\
        );

    \I__707\ : InMux
    port map (
            O => \N__7854\,
            I => \N__7841\
        );

    \I__706\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7841\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__7846\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7841\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__7836\,
            I => \N__7831\
        );

    \I__702\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7828\
        );

    \I__701\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7823\
        );

    \I__700\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7823\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__7828\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__7823\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__7818\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__7815\,
            I => \uu0.un4_l_count_16_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7809\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__7806\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__692\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7799\
        );

    \I__691\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7796\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__7799\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7796\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__688\ : IoInMux
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__7788\,
            I => \uu0.un11_l_count_i\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__7785\,
            I => \N__7782\
        );

    \I__685\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7776\
        );

    \I__684\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7773\
        );

    \I__683\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7768\
        );

    \I__682\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7768\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7765\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__7773\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__7768\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__7765\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__677\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__7755\,
            I => \uu0.un4_l_count_13\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__674\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7746\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__672\ : Span4Mux_s2_v
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__7740\,
            I => \uu2.mem0.N_139\
        );

    \I__670\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7731\
        );

    \I__668\ : IoSpan4Mux
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__7728\,
            I => \uart_RXD\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__665\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7716\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__7716\,
            I => \uu2.mem0.N_137\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__661\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__7704\,
            I => \uu2.mem0.N_141\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__7701\,
            I => \uu2.bitmap_pmux_u_0_a2_0_cascade_\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__656\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__7689\,
            I => \uu2.mem0.N_140\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__651\ : IoSpan4Mux
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__7677\,
            I => clk_in_c
        );

    \INVuu2.w_addr_user_7C\ : INV
    port map (
            O => \INVuu2.w_addr_user_7C_net\,
            I => \N__21656\
        );

    \INVuu2.w_addr_user_nesr_5C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_5C_net\,
            I => \N__21622\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__21645\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__21653\
        );

    \INVuu2.bitmap_168C\ : INV
    port map (
            O => \INVuu2.bitmap_168C_net\,
            I => \N__21659\
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__21649\
        );

    \INVuu2.w_addr_displaying_3_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_3_rep1C_net\,
            I => \N__21662\
        );

    \INVuu2.bitmap_194C\ : INV
    port map (
            O => \INVuu2.bitmap_194C_net\,
            I => \N__21669\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__21625\
        );

    \INVuu2.w_addr_user_nesr_8C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_8C_net\,
            I => \N__21648\
        );

    \INVuu2.w_addr_displaying_nesr_7C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_7C_net\,
            I => \N__21655\
        );

    \INVuu2.bitmap_186C\ : INV
    port map (
            O => \INVuu2.bitmap_186C_net\,
            I => \N__21661\
        );

    \INVuu2.w_addr_displaying_fast_2C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_2C_net\,
            I => \N__21668\
        );

    \INVuu2.w_addr_displaying_nesr_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_4C_net\,
            I => \N__21672\
        );

    \INVuu2.w_addr_user_4C\ : INV
    port map (
            O => \INVuu2.w_addr_user_4C_net\,
            I => \N__21654\
        );

    \INVuu2.w_addr_user_1C\ : INV
    port map (
            O => \INVuu2.w_addr_user_1C_net\,
            I => \N__21660\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9759\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \bu_rx_data_rdy_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19437\,
            GLOBALBUFFEROUTPUT => bu_rx_data_rdy_0_g
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11844\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7791\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15585\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__10329\,
            in1 => \N__11257\,
            in2 => \N__12927\,
            in3 => \N__9399\,
            lcout => \uu2.mem0.N_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__10330\,
            in1 => \N__12381\,
            in2 => \N__9585\,
            in3 => \N__11259\,
            lcout => \uu2.mem0.N_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIFPHP1_3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001000"
        )
    port map (
            in0 => \N__10706\,
            in1 => \N__9411\,
            in2 => \N__10604\,
            in3 => \N__10402\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_u_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIUI3J3_3_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110000"
        )
    port map (
            in0 => \N__10403\,
            in1 => \N__10600\,
            in2 => \N__7701\,
            in3 => \N__8109\,
            lcout => \uu2.N_922_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__10404\,
            in1 => \N__10331\,
            in2 => \N__9637\,
            in3 => \N__11258\,
            lcout => \uu2.mem0.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__11256\,
            in1 => \N__9858\,
            in2 => \N__10710\,
            in3 => \N__10328\,
            lcout => \uu2.mem0.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011110000"
        )
    port map (
            in0 => \N__9584\,
            in1 => \N__14084\,
            in2 => \N__9631\,
            in3 => \N__13997\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__19166\
        );

    \uu0.l_count_6_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__8809\,
            in2 => \N__9123\,
            in3 => \N__9084\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21646\,
            ce => \N__8725\,
            sr => \N__19216\
        );

    \buart.Z_rx.hh_1_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11558\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \buart.Z_rx.hh_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7737\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.l_precount_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.delay_line_1_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7803\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.delay_line_0_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7779\,
            in1 => \N__7835\,
            in2 => \N__7922\,
            in3 => \N__7855\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.l_precount_2_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7857\,
            in1 => \N__7917\,
            in2 => \_gnd_net_\,
            in3 => \N__7780\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.l_precount_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7916\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21641\,
            ce => 'H',
            sr => \N__19217\
        );

    \uu0.l_precount_3_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7781\,
            in1 => \N__7834\,
            in2 => \N__7923\,
            in3 => \N__7854\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21632\,
            ce => 'H',
            sr => \N__19218\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7853\,
            in1 => \N__8133\,
            in2 => \N__7836\,
            in3 => \N__7964\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI96A32_18_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8205\,
            in1 => \N__8741\,
            in2 => \N__7818\,
            in3 => \N__9085\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_11_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7758\,
            in1 => \N__8625\,
            in2 => \N__7815\,
            in3 => \N__7884\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_RNILLLG7_1_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7812\,
            in2 => \N__7806\,
            in3 => \N__7802\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2CNU_11_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__7873\,
            in2 => \N__7785\,
            in3 => \N__7984\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__7939\,
            in2 => \N__7992\,
            in3 => \N__7965\,
            lcout => \uu0.un66_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__7968\,
            in1 => \_gnd_net_\,
            in2 => \N__7947\,
            in3 => \N__7991\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__8726\,
            sr => \N__19220\
        );

    \uu0.l_count_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8803\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__8726\,
            sr => \N__19220\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7966\,
            in1 => \_gnd_net_\,
            in2 => \N__7946\,
            in3 => \N__7988\,
            lcout => OPEN,
            ltout => \uu0.un55_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_3_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__8640\,
            in1 => \_gnd_net_\,
            in2 => \N__7995\,
            in3 => \N__8805\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__8726\,
            sr => \N__19220\
        );

    \uu0.l_count_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7990\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__8726\,
            sr => \N__19220\
        );

    \uu0.l_count_11_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__7874\,
            in1 => \N__8073\,
            in2 => \N__8899\,
            in3 => \N__8804\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__8726\,
            sr => \N__19220\
        );

    \uu0.l_count_RNI04591_10_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8088\,
            in1 => \N__8059\,
            in2 => \N__8184\,
            in3 => \N__7938\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2GS72_4_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7921\,
            in1 => \N__8159\,
            in2 => \N__7887\,
            in3 => \N__8008\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__7875\,
            in2 => \N__8702\,
            in3 => \N__8060\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8183\,
            in1 => \N__8883\,
            in2 => \N__7860\,
            in3 => \N__8009\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => \N__8727\,
            sr => \N__19222\
        );

    \uu0.l_count_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8063\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => \N__8727\,
            sr => \N__19222\
        );

    \uu0.l_count_10_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8062\,
            in1 => \N__8700\,
            in2 => \N__8094\,
            in3 => \N__8885\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => \N__8727\,
            sr => \N__19222\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__8090\,
            in1 => \_gnd_net_\,
            in2 => \N__8703\,
            in3 => \N__8061\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_9_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8064\,
            in1 => \N__8884\,
            in2 => \_gnd_net_\,
            in3 => \N__8701\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => \N__8727\,
            sr => \N__19222\
        );

    \uu0.l_count_13_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__8031\,
            in1 => \N__8813\,
            in2 => \N__8040\,
            in3 => \N__8909\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21611\,
            ce => \N__8729\,
            sr => \N__19226\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8182\,
            in1 => \N__8221\,
            in2 => \_gnd_net_\,
            in3 => \N__8010\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8910\,
            in1 => \N__8814\,
            in2 => \N__8043\,
            in3 => \N__8204\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21611\,
            ce => \N__8729\,
            sr => \N__19226\
        );

    \uu0.l_count_12_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__8908\,
            in1 => \N__8022\,
            in2 => \N__8817\,
            in3 => \N__8222\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21611\,
            ce => \N__8729\,
            sr => \N__19226\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__8021\,
            in1 => \_gnd_net_\,
            in2 => \N__8223\,
            in3 => \_gnd_net_\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIFAQ9_13_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8030\,
            in2 => \_gnd_net_\,
            in3 => \N__8020\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => \uu0.un4_l_count_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8217\,
            in1 => \N__8203\,
            in2 => \N__8187\,
            in3 => \N__8181\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_4_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8949\,
            in1 => \N__8815\,
            in2 => \_gnd_net_\,
            in3 => \N__8157\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21611\,
            ce => \N__8729\,
            sr => \N__19226\
        );

    \uu0.l_count_5_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8950\,
            in1 => \N__8158\,
            in2 => \_gnd_net_\,
            in3 => \N__8132\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21604\,
            ce => \N__8730\,
            sr => \N__19229\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8160\,
            in2 => \_gnd_net_\,
            in3 => \N__8131\,
            lcout => \uu0.un88_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_2_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__12377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10400\,
            lcout => \uu2.N_34\,
            ltout => \uu2.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_5_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10700\,
            in1 => \N__10595\,
            in2 => \N__8112\,
            in3 => \N__9398\,
            lcout => \uu2.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIDKOL_0_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10399\,
            lcout => \uu2.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIV1P31_4_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__10699\,
            in1 => \N__12375\,
            in2 => \_gnd_net_\,
            in3 => \N__9397\,
            lcout => \uu2.N_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__10401\,
            in1 => \N__9042\,
            in2 => \N__12735\,
            in3 => \N__9716\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__9040\,
            in1 => \N__9709\,
            in2 => \N__11166\,
            in3 => \N__8253\,
            lcout => \uu2.mem0.N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__11255\,
            in1 => \N__9038\,
            in2 => \N__10335\,
            in3 => \N__10435\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__9714\,
            in1 => \N__13266\,
            in2 => \N__8289\,
            in3 => \N__8268\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__9710\,
            in1 => \N__9039\,
            in2 => \N__11331\,
            in3 => \N__10436\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIPAN5U_3_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__8274\,
            in1 => \N__10857\,
            in2 => \N__9423\,
            in3 => \N__10719\,
            lcout => \uu2.bitmap_pmux\,
            ltout => \uu2.bitmap_pmux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__8235\,
            in1 => \N__12783\,
            in2 => \N__8262\,
            in3 => \N__9715\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__9037\,
            in1 => \N__10324\,
            in2 => \N__8252\,
            in3 => \N__11254\,
            lcout => \uu2.mem0.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__11283\,
            in1 => \N__10437\,
            in2 => \N__9717\,
            in3 => \N__9041\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8569\,
            in1 => \N__8322\,
            in2 => \N__8356\,
            in3 => \N__8611\,
            lcout => \uu2.un404_ci\,
            ltout => \uu2.un404_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8421\,
            in1 => \N__8432\,
            in2 => \N__8439\,
            in3 => \N__8391\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21665\,
            ce => \N__8334\,
            sr => \N__19202\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8464\,
            in2 => \_gnd_net_\,
            in3 => \N__8532\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_7_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8380\,
            in1 => \N__8408\,
            in2 => \N__8415\,
            in3 => \N__8497\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21665\,
            ce => \N__8334\,
            sr => \N__19202\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8407\,
            in2 => \_gnd_net_\,
            in3 => \N__8379\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8533\,
            in1 => \N__8381\,
            in2 => \N__8471\,
            in3 => \N__8496\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21665\,
            ce => \N__8334\,
            sr => \N__19202\
        );

    \uu2.r_addr_esr_3_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8570\,
            in1 => \N__8323\,
            in2 => \N__8357\,
            in3 => \N__8612\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21665\,
            ce => \N__8334\,
            sr => \N__19202\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10121\,
            in2 => \_gnd_net_\,
            in3 => \N__19284\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_4_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000110101010"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__14076\,
            in2 => \N__12885\,
            in3 => \N__13990\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_4C_net\,
            ce => 'H',
            sr => \N__19167\
        );

    \uu2.r_addr_2_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10114\,
            in1 => \N__8607\,
            in2 => \N__8324\,
            in3 => \N__8565\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21647\,
            ce => 'H',
            sr => \N__19200\
        );

    \uu2.r_addr_4_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8525\,
            in1 => \N__8498\,
            in2 => \_gnd_net_\,
            in3 => \N__10115\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21647\,
            ce => 'H',
            sr => \N__19200\
        );

    \uu0.sec_clk_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13915\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21647\,
            ce => 'H',
            sr => \N__19200\
        );

    \uu2.r_addr_0_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8605\,
            in2 => \_gnd_net_\,
            in3 => \N__10116\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21642\,
            ce => 'H',
            sr => \N__19199\
        );

    \uu2.r_addr_1_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8564\,
            in1 => \N__8606\,
            in2 => \_gnd_net_\,
            in3 => \N__10117\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21642\,
            ce => 'H',
            sr => \N__19199\
        );

    \uu0.l_count_7_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8952\,
            in1 => \N__8802\,
            in2 => \N__9057\,
            in3 => \N__8674\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21633\,
            ce => \N__8724\,
            sr => \N__19219\
        );

    \uu2.r_addr_5_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8534\,
            in1 => \N__8499\,
            in2 => \N__10122\,
            in3 => \N__8460\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu2.trig_rd_det_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13860\,
            in2 => \_gnd_net_\,
            in3 => \N__10898\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu2.trig_rd_det_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10136\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu2.vram_rd_clk_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13861\,
            in2 => \_gnd_net_\,
            in3 => \N__8997\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu2.l_count_5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10027\,
            in1 => \N__10061\,
            in2 => \_gnd_net_\,
            in3 => \N__9269\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu2.l_count_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__9268\,
            in1 => \N__10003\,
            in2 => \_gnd_net_\,
            in3 => \N__9221\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__19201\
        );

    \uu0.l_count_17_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8835\,
            in1 => \N__8889\,
            in2 => \N__8658\,
            in3 => \N__8853\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21617\,
            ce => \N__8728\,
            sr => \N__19223\
        );

    \uu0.l_count_16_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8852\,
            in1 => \N__8801\,
            in2 => \N__8898\,
            in3 => \N__8834\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21617\,
            ce => \N__8728\,
            sr => \N__19223\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8936\,
            in1 => \N__9086\,
            in2 => \N__9122\,
            in3 => \N__8676\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__8653\,
            in2 => \N__8838\,
            in3 => \N__8833\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8800\,
            in2 => \N__8745\,
            in3 => \N__8742\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21617\,
            ce => \N__8728\,
            sr => \N__19223\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8693\,
            in1 => \N__8675\,
            in2 => \N__8657\,
            in3 => \N__8638\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9338\,
            in1 => \N__9006\,
            in2 => \N__9186\,
            in3 => \N__8958\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_9_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9223\,
            in1 => \N__10050\,
            in2 => \N__8978\,
            in3 => \N__9314\,
            lcout => OPEN,
            ltout => \uu2.un1_l_count_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9184\,
            in1 => \N__9342\,
            in2 => \N__9012\,
            in3 => \N__9005\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9267\,
            in2 => \N__9009\,
            in3 => \N__10051\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21612\,
            ce => 'H',
            sr => \N__19227\
        );

    \uu2.l_count_RNIFGGK1_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9241\,
            in1 => \N__10028\,
            in2 => \N__9144\,
            in3 => \N__9286\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__8996\,
            in1 => \N__9143\,
            in2 => \N__8979\,
            in3 => \N__9156\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21612\,
            ce => 'H',
            sr => \N__19227\
        );

    \uu2.l_count_3_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__9185\,
            in1 => \N__8995\,
            in2 => \N__9294\,
            in3 => \N__9198\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21612\,
            ce => 'H',
            sr => \N__19227\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9222\,
            in1 => \N__10049\,
            in2 => \N__8977\,
            in3 => \N__9313\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_7_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10005\,
            in1 => \N__9243\,
            in2 => \N__9270\,
            in3 => \N__9225\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21605\,
            ce => 'H',
            sr => \N__19230\
        );

    \uu2.l_count_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9318\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21605\,
            ce => 'H',
            sr => \N__19230\
        );

    \uu2.l_count_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21605\,
            ce => 'H',
            sr => \N__19230\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9316\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9339\,
            in1 => \N__9315\,
            in2 => \N__9293\,
            in3 => \N__9179\,
            lcout => \uu2.un306_ci\,
            ltout => \uu2.un306_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10004\,
            in1 => \N__9242\,
            in2 => \N__9228\,
            in3 => \N__9224\,
            lcout => \uu2.un350_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9197\,
            in2 => \_gnd_net_\,
            in3 => \N__9180\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21599\,
            ce => 'H',
            sr => \N__19232\
        );

    \uu2.l_count_8_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9139\,
            in2 => \_gnd_net_\,
            in3 => \N__9155\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21599\,
            ce => 'H',
            sr => \N__19232\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9109\,
            in2 => \_gnd_net_\,
            in3 => \N__9090\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIJQOL_2_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10831\,
            lcout => OPEN,
            ltout => \uu2.w_data_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI37MM2_3_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9380\,
            in1 => \N__10573\,
            in2 => \N__9045\,
            in3 => \N__10876\,
            lcout => \uu2.w_data_0_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_4_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__10686\,
            in1 => \N__10586\,
            in2 => \N__10653\,
            in3 => \N__9381\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_4C_net\,
            ce => \N__9515\,
            sr => \N__19174\
        );

    \uu2.w_addr_displaying_nesr_RNI7MSO_4_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12358\,
            in2 => \_gnd_net_\,
            in3 => \N__9376\,
            lcout => \uu2.bitmap_pmux_u_0_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIPFLE1_3_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001010000000"
        )
    port map (
            in0 => \N__10379\,
            in1 => \N__10572\,
            in2 => \N__9388\,
            in3 => \N__10684\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIDKOL_0_0_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12359\,
            in2 => \_gnd_net_\,
            in3 => \N__10378\,
            lcout => \uu2.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_RNIC9NT_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10374\,
            in1 => \N__12252\,
            in2 => \_gnd_net_\,
            in3 => \N__12183\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI4GV31_2_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110011010"
        )
    port map (
            in0 => \N__9474\,
            in1 => \N__9375\,
            in2 => \N__12263\,
            in3 => \N__10377\,
            lcout => \uu2.N_112_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI7JV31_2_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001110"
        )
    port map (
            in0 => \N__10376\,
            in1 => \N__12253\,
            in2 => \N__12579\,
            in3 => \N__9475\,
            lcout => \uu2.bitmap_pmux_sn_N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIGD5V_2_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001111111"
        )
    port map (
            in0 => \N__10380\,
            in1 => \N__12486\,
            in2 => \N__9477\,
            in3 => \N__9374\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_RNIT30I1_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12257\,
            in2 => \N__9345\,
            in3 => \N__12360\,
            lcout => \uu2.N_921_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_2_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__9476\,
            in1 => \N__10636\,
            in2 => \_gnd_net_\,
            in3 => \N__10476\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_2C_net\,
            ce => 'H',
            sr => \N__19173\
        );

    \uu2.w_addr_displaying_fast_RNI245H_2_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__10375\,
            in1 => \N__12091\,
            in2 => \_gnd_net_\,
            in3 => \N__9470\,
            lcout => \uu2.bitmap_pmux_sn_N_54_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__11100\,
            in1 => \N__11130\,
            in2 => \N__11062\,
            in3 => \N__12666\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__19171\
        );

    \uu2.bitmap_RNIBG4K_58_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9456\,
            in1 => \N__9450\,
            in2 => \_gnd_net_\,
            in3 => \N__10970\,
            lcout => \uu2.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_58_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__11102\,
            in1 => \N__11132\,
            in2 => \N__11064\,
            in3 => \N__12668\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__19171\
        );

    \uu2.bitmap_93_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__12669\,
            in1 => \N__11060\,
            in2 => \N__11136\,
            in3 => \N__11103\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__19171\
        );

    \uu2.bitmap_221_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__11101\,
            in1 => \N__11131\,
            in2 => \N__11063\,
            in3 => \N__12667\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__19171\
        );

    \uu2.bitmap_RNIRETJ1_93_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__12362\,
            in1 => \N__9444\,
            in2 => \N__9438\,
            in3 => \N__10986\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNIRETJ1Z0Z_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIHPJ64_3_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__10212\,
            in1 => \N__10579\,
            in2 => \N__9429\,
            in3 => \N__10426\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_27_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIIU8Q8_72_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10427\,
            in1 => \N__12318\,
            in2 => \N__9426\,
            in3 => \N__10884\,
            lcout => \uu2.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__10316\,
            in1 => \N__10789\,
            in2 => \N__12966\,
            in3 => \N__11250\,
            lcout => \uu2.mem0.N_135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__11251\,
            in1 => \N__10317\,
            in2 => \N__13962\,
            in3 => \N__12558\,
            lcout => \uu2.mem0.N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_7_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__12560\,
            in1 => \N__10793\,
            in2 => \N__10527\,
            in3 => \N__10847\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_7C_net\,
            ce => \N__9516\,
            sr => \N__19169\
        );

    \uu2.w_addr_displaying_ness_6_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011011110"
        )
    port map (
            in0 => \N__10848\,
            in1 => \N__10878\,
            in2 => \N__10800\,
            in3 => \N__10524\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_7C_net\,
            ce => \N__9516\,
            sr => \N__19169\
        );

    \uu2.w_addr_displaying_fast_nesr_7_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__10797\,
            in1 => \N__10846\,
            in2 => \N__10526\,
            in3 => \N__10980\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_7C_net\,
            ce => \N__9516\,
            sr => \N__19169\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_8_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__10845\,
            in1 => \N__10517\,
            in2 => \N__10799\,
            in3 => \N__12559\,
            lcout => \uu2.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0ES07_5_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__10844\,
            in2 => \N__10525\,
            in3 => \N__9685\,
            lcout => \uu2.w_addr_displaying_RNI0ES07Z0Z_5\,
            ltout => \uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI47N27_5_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9519\,
            in3 => \N__15584\,
            lcout => \uu2.N_32_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__12200\,
            in1 => \N__9661\,
            in2 => \N__10333\,
            in3 => \N__11252\,
            lcout => \uu2.mem0.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI20V6_8_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13954\,
            in1 => \N__9632\,
            in2 => \N__9663\,
            in3 => \N__9564\,
            lcout => \uu2.w_addr_user_3_i_a2_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100110"
        )
    port map (
            in0 => \N__9662\,
            in1 => \N__13955\,
            in2 => \N__14030\,
            in3 => \N__14063\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12815\,
            sr => \N__19168\
        );

    \uu2.w_addr_user_nesr_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__14060\,
            in1 => \N__9636\,
            in2 => \N__9857\,
            in3 => \N__9566\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12815\,
            sr => \N__19168\
        );

    \uu2.w_addr_user_nesr_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__9567\,
            in1 => \N__9815\,
            in2 => \N__12971\,
            in3 => \N__14059\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12815\,
            sr => \N__19168\
        );

    \uu2.w_addr_user_nesr_6_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__14062\,
            in1 => \N__14023\,
            in2 => \N__9870\,
            in3 => \N__9816\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12815\,
            sr => \N__19168\
        );

    \uu2.w_addr_user_nesr_RNO_0_3_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__9565\,
            in1 => \N__9798\,
            in2 => \N__9639\,
            in3 => \N__9850\,
            lcout => OPEN,
            ltout => \uu2.N_161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__14061\,
            in1 => \_gnd_net_\,
            in2 => \N__9645\,
            in3 => \N__12873\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12815\,
            sr => \N__19168\
        );

    \uu2.un28_w_addr_user_i_0_o2_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__11276\,
            in1 => \N__11007\,
            in2 => \N__11019\,
            in3 => \N__11206\,
            lcout => \uu2.N_101\,
            ltout => \uu2.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIE43C7_6_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__12967\,
            in1 => \N__9814\,
            in2 => \N__9642\,
            in3 => \N__10275\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIFBD5_3_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__9797\,
            in1 => \N__9846\,
            in2 => \N__9638\,
            in3 => \N__9574\,
            lcout => \uu2.N_106\,
            ltout => \uu2.N_106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNO_0_6_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__12962\,
            in1 => \N__12849\,
            in2 => \N__9873\,
            in3 => \N__12912\,
            lcout => \uu2.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNINJD5_3_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12911\,
            in1 => \N__9795\,
            in2 => \N__12852\,
            in3 => \N__9845\,
            lcout => OPEN,
            ltout => \uu2.w_addr_user_3_i_a2_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIPJCC_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9825\,
            in2 => \N__9819\,
            in3 => \_gnd_net_\,
            lcout => \uu2.N_230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__11207\,
            in1 => \N__9796\,
            in2 => \N__10334\,
            in3 => \N__10605\,
            lcout => \uu2.mem0.N_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12691\,
            in2 => \_gnd_net_\,
            in3 => \N__13916\,
            lcout => \oneSecStrb\,
            ltout => \oneSecStrb_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13090\,
            in1 => \N__14362\,
            in2 => \N__9762\,
            in3 => \N__14480\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21634\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__9758\,
            in1 => \N__10274\,
            in2 => \_gnd_net_\,
            in3 => \N__11204\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13917\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0_sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21634\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_i_o2_0_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10273\,
            in2 => \_gnd_net_\,
            in3 => \N__11203\,
            lcout => \uu2.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10297\,
            in1 => \N__11304\,
            in2 => \_gnd_net_\,
            in3 => \N__11205\,
            lcout => \uu2.mem0.N_54_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9969\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9957\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9945\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9933\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9921\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9909\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9897\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9885\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__11343\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111001110"
        )
    port map (
            in0 => \N__11543\,
            in1 => \N__13217\,
            in2 => \N__11523\,
            in3 => \N__11480\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \N__19224\
        );

    \buart.Z_tx.bitcount_0_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13216\,
            in1 => \N__11519\,
            in2 => \_gnd_net_\,
            in3 => \N__11542\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \N__19224\
        );

    \buart.Z_tx.bitcount_3_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__11544\,
            in1 => \N__11580\,
            in2 => \N__13218\,
            in3 => \N__11457\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \N__19224\
        );

    \buart.Z_tx.bitcount_2_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13212\,
            in2 => \_gnd_net_\,
            in3 => \N__11586\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \N__19224\
        );

    \buart.Z_rx.bitcount_es_1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__10182\,
            in1 => \N__12053\,
            in2 => \N__11685\,
            in3 => \N__11820\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21613\,
            ce => \N__12025\,
            sr => \N__19228\
        );

    \buart.Z_rx.bitcount_es_2_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__11819\,
            in1 => \N__10173\,
            in2 => \N__12060\,
            in3 => \N__11628\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21613\,
            ce => \N__12025\,
            sr => \N__19228\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10146\,
            in2 => \_gnd_net_\,
            in3 => \N__10137\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10029\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11867\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11681\,
            in2 => \_gnd_net_\,
            in3 => \N__10176\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11627\,
            in2 => \_gnd_net_\,
            in3 => \N__10167\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11711\,
            in2 => \_gnd_net_\,
            in3 => \N__10164\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__12057\,
            in1 => \N__11827\,
            in2 => \N__11655\,
            in3 => \N__10161\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21606\,
            ce => \N__12030\,
            sr => \N__19231\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11940\,
            in2 => \N__11772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11921\,
            in2 => \_gnd_net_\,
            in3 => \N__10158\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11821\,
            in1 => \N__11970\,
            in2 => \_gnd_net_\,
            in3 => \N__10155\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__21600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11987\,
            in2 => \_gnd_net_\,
            in3 => \N__10152\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__11823\,
            in1 => \N__11898\,
            in2 => \N__11958\,
            in3 => \N__10149\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__11822\,
            in1 => \N__10227\,
            in2 => \N__11925\,
            in3 => \N__11899\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_194_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__12437\,
            in1 => \N__13670\,
            in2 => \N__13420\,
            in3 => \N__13634\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.bitmap_RNII0BN_69_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100100111011"
        )
    port map (
            in0 => \N__12479\,
            in1 => \N__10979\,
            in2 => \N__10203\,
            in3 => \N__10188\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_25_i_m2_am_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIG91I1_66_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101100"
        )
    port map (
            in0 => \N__10221\,
            in1 => \N__10194\,
            in2 => \N__10215\,
            in3 => \N__12361\,
            lcout => \uu2.bitmap_RNIG91I1Z0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_34_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101101101"
        )
    port map (
            in0 => \N__13636\,
            in1 => \N__13414\,
            in2 => \N__13679\,
            in3 => \N__12439\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.bitmap_69_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101100110111"
        )
    port map (
            in0 => \N__12441\,
            in1 => \N__13678\,
            in2 => \N__13422\,
            in3 => \N__13638\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.bitmap_66_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000111101"
        )
    port map (
            in0 => \N__13637\,
            in1 => \N__13415\,
            in2 => \N__13680\,
            in3 => \N__12440\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.bitmap_197_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__12438\,
            in1 => \N__13671\,
            in2 => \N__13421\,
            in3 => \N__13635\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.w_addr_displaying_fast_0_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__10485\,
            in1 => \_gnd_net_\,
            in2 => \N__12488\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__19177\
        );

    \uu2.w_addr_displaying_3_rep1_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__10695\,
            in1 => \N__10483\,
            in2 => \N__10648\,
            in3 => \N__12262\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_2_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__10479\,
            in1 => \N__10637\,
            in2 => \_gnd_net_\,
            in3 => \N__10697\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_fast_3_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__10696\,
            in1 => \N__10484\,
            in2 => \N__10649\,
            in3 => \N__12095\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__10482\,
            in1 => \N__10698\,
            in2 => \N__10596\,
            in3 => \N__10638\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_0_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10477\,
            in2 => \_gnd_net_\,
            in3 => \N__12374\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_8_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__10481\,
            in1 => \N__10539\,
            in2 => \_gnd_net_\,
            in3 => \N__12195\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_5_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__10513\,
            in1 => \N__10480\,
            in2 => \_gnd_net_\,
            in3 => \N__10843\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.w_addr_displaying_1_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__10478\,
            in1 => \N__10425\,
            in2 => \_gnd_net_\,
            in3 => \N__10391\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__19175\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__10332\,
            in1 => \N__10830\,
            in2 => \N__11253\,
            in3 => \N__12850\,
            lcout => \uu2.mem0.N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIFJI02_212_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111100"
        )
    port map (
            in0 => \N__13689\,
            in1 => \N__12547\,
            in2 => \N__13791\,
            in3 => \N__12447\,
            lcout => \uu2.bitmap_RNIFJI02Z0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNI6J081_6_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12191\,
            in1 => \_gnd_net_\,
            in2 => \N__12567\,
            in3 => \N__10783\,
            lcout => \uu2.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNI12TI1_0_6_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__10788\,
            in2 => \N__12581\,
            in3 => \N__12194\,
            lcout => \uu2.bitmap_pmux_u_0_83_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNI12TI1_1_6_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001000010"
        )
    port map (
            in0 => \N__12192\,
            in1 => \N__12571\,
            in2 => \N__10798\,
            in3 => \N__10828\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNI12TI1_6_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101110111"
        )
    port map (
            in0 => \N__10827\,
            in1 => \N__10787\,
            in2 => \N__12582\,
            in3 => \N__12193\,
            lcout => OPEN,
            ltout => \uu2.N_100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI3OPR5_2_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__10752\,
            in1 => \N__10746\,
            in2 => \N__10740\,
            in3 => \N__10737\,
            lcout => OPEN,
            ltout => \uu2.N_923_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8ND5G_3_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__10731\,
            in1 => \N__10932\,
            in2 => \N__10722\,
            in3 => \N__12279\,
            lcout => \uu2.w_addr_displaying_RNI8ND5GZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_314_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100111"
        )
    port map (
            in0 => \N__11119\,
            in1 => \N__11049\,
            in2 => \N__11089\,
            in3 => \N__12652\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__19172\
        );

    \uu2.bitmap_218_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__12651\,
            in1 => \N__11079\,
            in2 => \N__11061\,
            in3 => \N__11118\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__19172\
        );

    \uu2.bitmap_90_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000110101"
        )
    port map (
            in0 => \N__11120\,
            in1 => \N__11050\,
            in2 => \N__11090\,
            in3 => \N__12653\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__19172\
        );

    \uu2.bitmap_RNI6H8O_90_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__10978\,
            in1 => \N__12489\,
            in2 => \N__11001\,
            in3 => \N__10992\,
            lcout => \uu2.bitmap_pmux_25_i_m2_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIU0UJ_314_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__12096\,
            in1 => \N__10977\,
            in2 => \_gnd_net_\,
            in3 => \N__10925\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_21_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIBNS22_180_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000001110"
        )
    port map (
            in0 => \N__13806\,
            in1 => \N__12264\,
            in2 => \N__10950\,
            in3 => \N__12135\,
            lcout => OPEN,
            ltout => \uu2.N_393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_RNIN52C4_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10947\,
            in2 => \N__10935\,
            in3 => \N__10911\,
            lcout => \uu2.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI05EB1_314_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10926\,
            in1 => \N__12199\,
            in2 => \_gnd_net_\,
            in3 => \N__10917\,
            lcout => \uu2.N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__13875\,
            in1 => \N__10905\,
            in2 => \N__13199\,
            in3 => \N__19287\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIITTD7_6_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15574\,
            in2 => \_gnd_net_\,
            in3 => \N__13980\,
            lcout => \uu2.un28_w_addr_user_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__18006\,
            in1 => \N__18046\,
            in2 => \_gnd_net_\,
            in3 => \N__19949\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__18047\,
            in1 => \N__15810\,
            in2 => \N__11139\,
            in3 => \N__15843\,
            lcout => \Lab_UT.didp.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIFKHR3_1_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17964\,
            in1 => \N__14571\,
            in2 => \_gnd_net_\,
            in3 => \N__17319\,
            lcout => \Lab_UT.sec2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIHMHR3_2_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14570\,
            in1 => \N__16044\,
            in2 => \_gnd_net_\,
            in3 => \N__17295\,
            lcout => \Lab_UT.sec2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIJOHR3_3_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15999\,
            in1 => \N__14572\,
            in2 => \_gnd_net_\,
            in3 => \N__17265\,
            lcout => \Lab_UT.sec2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_a2_0_4_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11303\,
            in1 => \N__11156\,
            in2 => \N__12779\,
            in3 => \N__11321\,
            lcout => \uu2.un28_w_addr_user_i_0_a2_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13079\,
            in1 => \N__14356\,
            in2 => \_gnd_net_\,
            in3 => \N__14483\,
            lcout => \Lab_UT.dispString.un42_dOutP\,
            ltout => \Lab_UT.dispString.un42_dOutP_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__11355\,
            in1 => \N__11349\,
            in2 => \N__11010\,
            in3 => \N__12636\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_a2_0_0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12721\,
            in2 => \_gnd_net_\,
            in3 => \N__13256\,
            lcout => \uu2.un28_w_addr_user_i_0_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111010101"
        )
    port map (
            in0 => \N__14481\,
            in1 => \N__17577\,
            in2 => \N__14366\,
            in3 => \N__17436\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010111010"
        )
    port map (
            in0 => \N__13080\,
            in1 => \N__14357\,
            in2 => \N__11358\,
            in3 => \N__14482\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__12612\,
            in1 => \N__13084\,
            in2 => \_gnd_net_\,
            in3 => \N__12621\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__12411\,
            in1 => \N__11600\,
            in2 => \N__13091\,
            in3 => \N__17294\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001111"
        )
    port map (
            in0 => \N__14476\,
            in1 => \N__11601\,
            in2 => \N__13092\,
            in3 => \N__13239\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21626\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__13839\,
            in1 => \N__13821\,
            in2 => \_gnd_net_\,
            in3 => \N__19278\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__14253\,
            in1 => \N__14965\,
            in2 => \N__14488\,
            in3 => \N__16638\,
            lcout => \Lab_UT.dispString.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_0_a3_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11155\,
            in1 => \N__11320\,
            in2 => \N__12725\,
            in3 => \N__13255\,
            lcout => OPEN,
            ltout => \uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_0_a3_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12766\,
            in1 => \N__11302\,
            in2 => \N__11286\,
            in3 => \N__11275\,
            lcout => \uu2.un1_w_user_cr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101111110"
        )
    port map (
            in0 => \N__14365\,
            in1 => \N__13089\,
            in2 => \N__14489\,
            in3 => \N__12675\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21626\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__13183\,
            in1 => \N__11412\,
            in2 => \_gnd_net_\,
            in3 => \N__11451\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11445\,
            in2 => \_gnd_net_\,
            in3 => \N__13181\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.uart_tx_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__13182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11439\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_2_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11400\,
            in1 => \N__13184\,
            in2 => \_gnd_net_\,
            in3 => \N__11418\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__13185\,
            in1 => \N__11388\,
            in2 => \_gnd_net_\,
            in3 => \N__11406\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_4_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11376\,
            in1 => \N__13186\,
            in2 => \_gnd_net_\,
            in3 => \N__11394\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_5_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__13187\,
            in1 => \N__11364\,
            in2 => \_gnd_net_\,
            in3 => \N__11382\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.shifter_6_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13224\,
            in1 => \N__13188\,
            in2 => \_gnd_net_\,
            in3 => \N__11370\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => \N__13115\,
            sr => \N__19221\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__11475\,
            in1 => \N__11568\,
            in2 => \N__11498\,
            in3 => \N__13338\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11604\,
            in3 => \N__13180\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIFV4E_1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14297\,
            in2 => \_gnd_net_\,
            in3 => \N__14407\,
            lcout => \Lab_UT.dispString.N_191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100111001100"
        )
    port map (
            in0 => \N__11517\,
            in1 => \N__11494\,
            in2 => \N__11481\,
            in3 => \N__11540\,
            lcout => \buart.Z_tx.bitcount_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__11579\,
            in1 => \N__11516\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.uart_busy_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14653\,
            in1 => \N__11562\,
            in2 => \_gnd_net_\,
            in3 => \N__11745\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__11541\,
            in1 => \N__11518\,
            in2 => \N__11499\,
            in3 => \N__11479\,
            lcout => \buart.Z_tx.un1_bitcount_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__11796\,
            in2 => \N__11904\,
            in3 => \N__11744\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13009\,
            in2 => \_gnd_net_\,
            in3 => \N__12986\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12985\,
            in1 => \N__13364\,
            in2 => \N__13011\,
            in3 => \N__13272\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11743\,
            in2 => \_gnd_net_\,
            in3 => \N__18986\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21399\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13008\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11626\,
            in1 => \N__11651\,
            in2 => \N__11712\,
            in3 => \N__11679\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIQ0DP_4_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11650\,
            in2 => \_gnd_net_\,
            in3 => \N__11624\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11680\,
            in1 => \N__11706\,
            in2 => \N__11748\,
            in3 => \N__11865\,
            lcout => \buart.Z_rx.idle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__11707\,
            in1 => \N__12059\,
            in2 => \N__11724\,
            in3 => \N__11829\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21601\,
            ce => \N__12026\,
            sr => \N__19233\
        );

    \buart.Z_rx.bitcount_es_RNINTCP_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11705\,
            in2 => \_gnd_net_\,
            in3 => \N__11864\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11678\,
            in1 => \N__11649\,
            in2 => \N__11631\,
            in3 => \N__11625\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__11866\,
            in1 => \N__12058\,
            in2 => \N__15759\,
            in3 => \N__11828\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21601\,
            ce => \N__12026\,
            sr => \N__19233\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__11824\,
            in1 => \_gnd_net_\,
            in2 => \N__11771\,
            in3 => \N__11939\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__11900\,
            in1 => \N__11825\,
            in2 => \N__11991\,
            in3 => \N__11997\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11986\,
            in1 => \N__11969\,
            in2 => \N__11957\,
            in3 => \N__11938\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11920\,
            in2 => \N__11907\,
            in3 => \N__11763\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__11877\,
            in1 => \_gnd_net_\,
            in2 => \N__11871\,
            in3 => \N__11868\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11764\,
            in2 => \_gnd_net_\,
            in3 => \N__11826\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_5_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18875\,
            in1 => \N__20161\,
            in2 => \N__21355\,
            in3 => \N__19933\,
            lcout => \Lab_UT.dictrl.g1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIJAJ21_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18494\,
            in1 => \N__21348\,
            in2 => \N__20937\,
            in3 => \N__18876\,
            lcout => \Lab_UT.dictrl.g0_17_a6_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_168_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011001010110"
        )
    port map (
            in0 => \N__13437\,
            in1 => \N__13603\,
            in2 => \N__13547\,
            in3 => \N__13576\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__19180\
        );

    \uu2.bitmap_RNISSSN_162_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12108\,
            in1 => \N__12090\,
            in2 => \_gnd_net_\,
            in3 => \N__12129\,
            lcout => \uu2.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011100011111"
        )
    port map (
            in0 => \N__13439\,
            in1 => \N__13607\,
            in2 => \N__13548\,
            in3 => \N__13578\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__19180\
        );

    \uu2.bitmap_203_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__13577\,
            in1 => \N__13530\,
            in2 => \N__13608\,
            in3 => \N__13438\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__19180\
        );

    \uu2.bitmap_RNIM9P11_75_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011101010101"
        )
    port map (
            in0 => \N__12578\,
            in1 => \N__12123\,
            in2 => \N__12117\,
            in3 => \N__12475\,
            lcout => \uu2.bitmap_pmux_24_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000110110"
        )
    port map (
            in0 => \N__12435\,
            in1 => \N__13404\,
            in2 => \N__13658\,
            in3 => \N__13621\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__19180\
        );

    \uu2.bitmap_290_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100011001"
        )
    port map (
            in0 => \N__13622\,
            in1 => \N__13654\,
            in2 => \N__13419\,
            in3 => \N__12436\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__19180\
        );

    \uu2.bitmap_RNI4LQU_34_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__12102\,
            in1 => \N__12089\,
            in2 => \N__12201\,
            in3 => \N__12066\,
            lcout => \uu2.bitmap_pmux_15_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100111"
        )
    port map (
            in0 => \N__13600\,
            in1 => \N__13452\,
            in2 => \N__13549\,
            in3 => \N__13573\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__19178\
        );

    \uu2.bitmap_200_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__13572\,
            in1 => \N__13537\,
            in2 => \N__13455\,
            in3 => \N__13599\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__19178\
        );

    \uu2.bitmap_72_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000110101"
        )
    port map (
            in0 => \N__13602\,
            in1 => \N__13454\,
            in2 => \N__13551\,
            in3 => \N__13575\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__19178\
        );

    \uu2.bitmap_RNI5T9T1_72_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__12402\,
            in1 => \N__12396\,
            in2 => \N__12390\,
            in3 => \N__12373\,
            lcout => \uu2.bitmap_RNI5T9T1Z0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011011011101111"
        )
    port map (
            in0 => \N__13601\,
            in1 => \N__13453\,
            in2 => \N__13550\,
            in3 => \N__13574\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__19178\
        );

    \uu2.bitmap_RNIGQ8J1_111_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12306\,
            in1 => \N__13881\,
            in2 => \_gnd_net_\,
            in3 => \N__12297\,
            lcout => OPEN,
            ltout => \uu2.N_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIL9SE4_2_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12291\,
            in2 => \N__12282\,
            in3 => \N__12207\,
            lcout => \uu2.N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIURJN1_40_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__12270\,
            in1 => \N__12258\,
            in2 => \N__12225\,
            in3 => \N__12213\,
            lcout => \uu2.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011101"
        )
    port map (
            in0 => \N__13773\,
            in1 => \N__13746\,
            in2 => \N__14232\,
            in3 => \N__13716\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__19176\
        );

    \uu2.bitmap_RNIU2IS_52_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12588\,
            in1 => \N__12190\,
            in2 => \_gnd_net_\,
            in3 => \N__12141\,
            lcout => \uu2.bitmap_RNIU2ISZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_52_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__13774\,
            in1 => \N__13747\,
            in2 => \N__14233\,
            in3 => \N__13717\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__19176\
        );

    \uu2.bitmap_84_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__13775\,
            in1 => \N__13748\,
            in2 => \N__14234\,
            in3 => \N__13718\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__19176\
        );

    \uu2.bitmap_87_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__13776\,
            in1 => \N__13749\,
            in2 => \N__14235\,
            in3 => \N__13719\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__19176\
        );

    \uu2.bitmap_RNIG5UR_84_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__12580\,
            in1 => \N__12504\,
            in2 => \N__12498\,
            in3 => \N__12487\,
            lcout => \uu2.bitmap_pmux_24_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI8CKM3_1_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16823\,
            in1 => \N__14564\,
            in2 => \_gnd_net_\,
            in3 => \N__15386\,
            lcout => \Lab_UT.sec1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNIAEKM3_2_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14563\,
            in1 => \N__15633\,
            in2 => \_gnd_net_\,
            in3 => \N__17573\,
            lcout => \Lab_UT.sec1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNILUSP3_1_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14580\,
            in1 => \N__14125\,
            in2 => \_gnd_net_\,
            in3 => \N__14180\,
            lcout => \Lab_UT.min1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_1_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20303\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21638\,
            ce => \N__16604\,
            sr => \N__19209\
        );

    \Lab_UT.dispString.dOut_RNO_3_2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__12702\,
            in1 => \N__13928\,
            in2 => \_gnd_net_\,
            in3 => \N__14159\,
            lcout => \Lab_UT.dispString.un46_dOutP_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_2_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20766\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21638\,
            ce => \N__16604\,
            sr => \N__19209\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIH9JB1_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__15426\,
            in1 => \N__16843\,
            in2 => \N__12606\,
            in3 => \N__18034\,
            lcout => \Lab_UT.didp.did_alarmMatch_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIDIHR3_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12604\,
            in1 => \N__14561\,
            in2 => \_gnd_net_\,
            in3 => \N__18035\,
            lcout => \Lab_UT.sec2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI6AKM3_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__14562\,
            in1 => \_gnd_net_\,
            in2 => \N__15435\,
            in3 => \N__16844\,
            lcout => \Lab_UT.sec1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__12635\,
            in1 => \N__17768\,
            in2 => \N__19290\,
            in3 => \N__17834\,
            lcout => \G_190\,
            ltout => \G_190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010001110101"
        )
    port map (
            in0 => \N__14335\,
            in1 => \N__14456\,
            in2 => \N__12624\,
            in3 => \N__12605\,
            lcout => \Lab_UT.dispString.i21_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100110011"
        )
    port map (
            in0 => \N__17505\,
            in1 => \N__14334\,
            in2 => \N__16848\,
            in3 => \N__14471\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m28_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000001010"
        )
    port map (
            in0 => \N__14472\,
            in1 => \N__15011\,
            in2 => \N__12615\,
            in3 => \N__17172\,
            lcout => \Lab_UT.dispString.N_204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19955\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21629\,
            ce => \N__18663\,
            sr => \N__19206\
        );

    \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__12972\,
            in1 => \N__12842\,
            in2 => \N__12881\,
            in3 => \N__12925\,
            lcout => \uu2.N_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_5_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011010010"
        )
    port map (
            in0 => \N__12926\,
            in1 => \N__12877\,
            in2 => \N__12851\,
            in3 => \N__14077\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_5C_net\,
            ce => \N__12816\,
            sr => \N__19170\
        );

    \Lab_UT.dictrl.m59_ns_1_ns_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16203\,
            lcout => \Lab_UT.dictrl.m59_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_3_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15752\,
            in1 => \N__15774\,
            in2 => \N__12804\,
            in3 => \N__14625\,
            lcout => \G_193\,
            ltout => \G_193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__14340\,
            in1 => \N__14441\,
            in2 => \N__12795\,
            in3 => \N__17264\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__12792\,
            in1 => \_gnd_net_\,
            in2 => \N__12786\,
            in3 => \N__13069\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_6_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100010"
        )
    port map (
            in0 => \N__17769\,
            in1 => \N__15500\,
            in2 => \N__12753\,
            in3 => \N__17835\,
            lcout => \G_189\,
            ltout => \G_189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12744\,
            in3 => \N__12741\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_5_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110100"
        )
    port map (
            in0 => \N__12701\,
            in1 => \N__13918\,
            in2 => \N__14361\,
            in3 => \N__14615\,
            lcout => \Lab_UT.dispString.m44_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13506\,
            in1 => \N__13068\,
            in2 => \_gnd_net_\,
            in3 => \N__14496\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111110001"
        )
    port map (
            in0 => \N__14336\,
            in1 => \N__15005\,
            in2 => \N__13085\,
            in3 => \N__14614\,
            lcout => \Lab_UT.dispString.m42_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__13201\,
            in1 => \N__13125\,
            in2 => \_gnd_net_\,
            in3 => \N__13233\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21610\,
            ce => \N__13119\,
            sr => \N__19225\
        );

    \buart.Z_tx.shifter_8_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13200\,
            in2 => \_gnd_net_\,
            in3 => \N__13134\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21610\,
            ce => \N__13119\,
            sr => \N__19225\
        );

    \Lab_UT.dispString.cnt_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14455\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21603\,
            ce => 'H',
            sr => \N__19204\
        );

    \Lab_UT.dispString.cnt_0_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__14310\,
            in1 => \N__14454\,
            in2 => \N__13078\,
            in3 => \N__15012\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21603\,
            ce => 'H',
            sr => \N__19204\
        );

    \Lab_UT.dispString.cnt_2_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__14453\,
            in1 => \N__14312\,
            in2 => \_gnd_net_\,
            in3 => \N__13055\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21603\,
            ce => 'H',
            sr => \N__19204\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13010\,
            in2 => \N__12990\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13365\,
            in2 => \_gnd_net_\,
            in3 => \N__13353\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__21598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13340\,
            in1 => \N__13281\,
            in2 => \_gnd_net_\,
            in3 => \N__13350\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__21598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13308\,
            in3 => \N__13347\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__21598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__13341\,
            in1 => \_gnd_net_\,
            in2 => \N__13320\,
            in3 => \N__13344\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__21598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__13295\,
            in1 => \N__13339\,
            in2 => \_gnd_net_\,
            in3 => \N__13323\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13316\,
            in1 => \N__13304\,
            in2 => \N__13296\,
            in3 => \N__13280\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUJLP6_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001000"
        )
    port map (
            in0 => \N__16290\,
            in1 => \N__14844\,
            in2 => \N__21261\,
            in3 => \N__19641\,
            lcout => \Lab_UT.dictrl.N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14660\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21594\,
            ce => \N__19316\,
            sr => \N__19235\
        );

    \buart.Z_rx.shifter_fast_7_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21594\,
            ce => \N__19316\,
            sr => \N__19235\
        );

    \buart.Z_rx.shifter_fast_6_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20362\,
            lcout => \buart__rx_shifter_fast_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21594\,
            ce => \N__19316\,
            sr => \N__19235\
        );

    \buart.Z_rx.shifter_6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21594\,
            ce => \N__19316\,
            sr => \N__19235\
        );

    \Lab_UT.dictrl.state_0_esr_RNIU7683_2_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16449\,
            in1 => \N__20029\,
            in2 => \N__19810\,
            in3 => \N__13377\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI88DT7_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__19665\,
            in1 => \N__21250\,
            in2 => \N__13371\,
            in3 => \N__14877\,
            lcout => \Lab_UT.dictrl.N_90_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m30_0_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__14896\,
            in1 => \_gnd_net_\,
            in2 => \N__18429\,
            in3 => \N__18941\,
            lcout => \Lab_UT.dictrl.m30_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_17_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18424\,
            in1 => \N__16131\,
            in2 => \N__16519\,
            in3 => \N__18942\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_14_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16732\,
            in1 => \N__16448\,
            in2 => \N__13368\,
            in3 => \N__19497\,
            lcout => \Lab_UT.dictrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIHC6L_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__14734\,
            in1 => \N__16367\,
            in2 => \N__21044\,
            in3 => \N__20929\,
            lcout => \Lab_UT.dictrl.g0_17_a6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNINEHL_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__18868\,
            in1 => \N__16259\,
            in2 => \N__21104\,
            in3 => \N__18381\,
            lcout => \Lab_UT.dictrl.g0_17_a6_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_17_a6_1_6_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19496\,
            in1 => \N__20374\,
            in2 => \N__21356\,
            in3 => \N__20595\,
            lcout => \Lab_UT.dictrl.g0_17_a6_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNI7FC61_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16380\,
            in1 => \N__18753\,
            in2 => \N__20163\,
            in3 => \N__20934\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_17_a6_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIU4P66_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__13491\,
            in1 => \N__13485\,
            in2 => \N__13479\,
            in3 => \N__13467\,
            lcout => \Lab_UT.dictrl.g0_17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_17_o6_1_4_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19495\,
            in1 => \N__20142\,
            in2 => \N__18633\,
            in3 => \N__18380\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIG3243_1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13461\,
            in2 => \N__13476\,
            in3 => \N__13473\,
            lcout => \Lab_UT.dictrl.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIO3GC_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16710\,
            in2 => \_gnd_net_\,
            in3 => \N__16258\,
            lcout => \Lab_UT.dictrl.g0_17_a6_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_17_o6_1_5_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__18428\,
            in1 => \N__18867\,
            in2 => \N__16731\,
            in3 => \N__20594\,
            lcout => \Lab_UT.dictrl.g0_17_o6_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15062\,
            in1 => \N__17208\,
            in2 => \_gnd_net_\,
            in3 => \N__14135\,
            lcout => \Lab_UT.didp.countrce4.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNIEQ8R3_3_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14568\,
            in1 => \N__17088\,
            in2 => \_gnd_net_\,
            in3 => \N__17358\,
            lcout => \Lab_UT.min2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIP2TP3_3_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15476\,
            in1 => \N__14569\,
            in2 => \_gnd_net_\,
            in3 => \N__16634\,
            lcout => \Lab_UT.min1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIN0TP3_2_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14566\,
            in1 => \N__15061\,
            in2 => \_gnd_net_\,
            in3 => \N__14163\,
            lcout => \Lab_UT.min1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIJSSP3_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17171\,
            in1 => \N__17207\,
            in2 => \_gnd_net_\,
            in3 => \N__14567\,
            lcout => \Lab_UT.min1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__17203\,
            in1 => \N__15184\,
            in2 => \_gnd_net_\,
            in3 => \N__19948\,
            lcout => \Lab_UT.didp.countrce4.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_1_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__17051\,
            in1 => \N__20304\,
            in2 => \N__16953\,
            in3 => \N__17004\,
            lcout => \Lab_UT.didp.countrce3.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__17204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14136\,
            lcout => \Lab_UT.didp.reset_12_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNIAM8R3_1_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14583\,
            in1 => \N__17003\,
            in2 => \_gnd_net_\,
            in3 => \N__17465\,
            lcout => \Lab_UT.min2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNI8K8R3_0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17050\,
            in1 => \N__14582\,
            in2 => \_gnd_net_\,
            in3 => \N__17504\,
            lcout => \Lab_UT.min2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNICO8R3_2_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14581\,
            in1 => \N__16904\,
            in2 => \_gnd_net_\,
            in3 => \N__17435\,
            lcout => \Lab_UT.min2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101011111"
        )
    port map (
            in0 => \N__17466\,
            in1 => \N__15013\,
            in2 => \N__14490\,
            in3 => \N__14184\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100111"
        )
    port map (
            in0 => \N__14367\,
            in1 => \N__14487\,
            in2 => \N__13509\,
            in3 => \N__16824\,
            lcout => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_7_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000110101010"
        )
    port map (
            in0 => \N__13953\,
            in1 => \N__14085\,
            in2 => \N__14031\,
            in3 => \N__13998\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.bitmap_111_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13929\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.vram_rd_clk_det_0_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.vram_rd_clk_det_1_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13835\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.bitmap_180_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__13777\,
            in1 => \N__13750\,
            in2 => \N__14229\,
            in3 => \N__13720\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.bitmap_215_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__13722\,
            in1 => \N__13779\,
            in2 => \N__14231\,
            in3 => \N__13752\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \uu2.bitmap_212_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__13778\,
            in1 => \N__13751\,
            in2 => \N__14230\,
            in3 => \N__13721\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__19179\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__16941\,
            in1 => \N__17052\,
            in2 => \_gnd_net_\,
            in3 => \N__19929\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNICGKM3_3_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14565\,
            in1 => \N__15339\,
            in2 => \_gnd_net_\,
            in3 => \N__17543\,
            lcout => \Lab_UT.sec1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIAC7D1_1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__14179\,
            in1 => \N__15050\,
            in2 => \N__14134\,
            in3 => \N__14155\,
            lcout => \Lab_UT.didp.did_alarmMatch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__14132\,
            in1 => \N__20302\,
            in2 => \N__15196\,
            in3 => \N__17206\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__15097\,
            in1 => \N__15138\,
            in2 => \N__14139\,
            in3 => \N__14133\,
            lcout => \Lab_UT.didp.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14124\,
            in2 => \_gnd_net_\,
            in3 => \N__17205\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__15060\,
            in1 => \N__20765\,
            in2 => \N__14094\,
            in3 => \N__15188\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15051\,
            in1 => \N__15137\,
            in2 => \N__14091\,
            in3 => \N__15098\,
            lcout => \Lab_UT.didp.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100001100"
        )
    port map (
            in0 => \N__21260\,
            in1 => \N__14598\,
            in2 => \N__17853\,
            in3 => \N__19647\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__21100\,
            in2 => \N__14088\,
            in3 => \N__20924\,
            lcout => \Lab_UT.dictrl.state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21644\,
            ce => \N__15872\,
            sr => \N__19210\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNI036C1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__19418\,
            in1 => \N__18738\,
            in2 => \N__18477\,
            in3 => \N__19757\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIH9933_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20923\,
            in2 => \N__14586\,
            in3 => \N__14502\,
            lcout => \Lab_UT.i16_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNIRKP91_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__19417\,
            in1 => \N__19646\,
            in2 => \N__18258\,
            in3 => \N__14694\,
            lcout => \Lab_UT.dictrl.i18_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__14458\,
            in1 => \N__17318\,
            in2 => \N__14364\,
            in3 => \N__15704\,
            lcout => \Lab_UT.dispString.dOut_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20930\,
            in1 => \N__19649\,
            in2 => \N__21259\,
            in3 => \N__19774\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100101111"
        )
    port map (
            in0 => \N__14457\,
            in1 => \N__17544\,
            in2 => \N__14363\,
            in3 => \N__17357\,
            lcout => \Lab_UT.dispString.m49_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_2_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18060\,
            in2 => \_gnd_net_\,
            in3 => \N__17950\,
            lcout => \Lab_UT.didp.countrce1.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18061\,
            in1 => \N__16035\,
            in2 => \_gnd_net_\,
            in3 => \N__17951\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17998\,
            in1 => \N__20491\,
            in2 => \N__14241\,
            in3 => \N__15993\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__15806\,
            in1 => \N__15994\,
            in2 => \N__14238\,
            in3 => \N__15842\,
            lcout => \Lab_UT.didp.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_idle_1_0_iclk_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__15582\,
            in1 => \N__17761\,
            in2 => \_gnd_net_\,
            in3 => \N__17819\,
            lcout => \Lab_UT.un1_idle_1_0_iclkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21217\,
            in1 => \N__19648\,
            in2 => \N__17628\,
            in3 => \N__19743\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicAlarmTrig_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17762\,
            in2 => \_gnd_net_\,
            in3 => \N__17820\,
            lcout => \G_186\,
            ltout => \G_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_4_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__17763\,
            in1 => \N__19282\,
            in2 => \N__14619\,
            in3 => \N__14616\,
            lcout => \G_191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_10_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20167\,
            in2 => \_gnd_net_\,
            in3 => \N__20608\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__19744\,
            in1 => \N__19650\,
            in2 => \N__14601\,
            in3 => \N__20386\,
            lcout => \Lab_UT.dictrl.G_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNIRFD0E_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17901\,
            in1 => \N__16106\,
            in2 => \N__18175\,
            in3 => \N__16073\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__15918\,
            in1 => \N__19009\,
            in2 => \N__14589\,
            in3 => \N__14693\,
            lcout => \Lab_UT.dicRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21620\,
            ce => 'H',
            sr => \N__19203\
        );

    \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__19286\,
            in1 => \N__20886\,
            in2 => \N__21237\,
            in3 => \N__14691\,
            lcout => \Lab_UT.didp.regrce4.LdAMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14692\,
            in1 => \N__17634\,
            in2 => \N__15024\,
            in3 => \N__21204\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21620\,
            ce => 'H',
            sr => \N__19203\
        );

    \Lab_UT.didp.ce_RNI51AM_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14673\,
            in2 => \_gnd_net_\,
            in3 => \N__15927\,
            lcout => \Lab_UT.didp.un1_dicLdSones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15941\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21620\,
            ce => 'H',
            sr => \N__19203\
        );

    \Lab_UT.didp.ce_RNI5U3I_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14667\,
            in2 => \_gnd_net_\,
            in3 => \N__14748\,
            lcout => \Lab_UT.didp.un1_dicLdStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_rep1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14654\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21614\,
            ce => \N__19318\,
            sr => \N__19234\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__18720\,
            in1 => \_gnd_net_\,
            in2 => \N__16376\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16359\,
            in2 => \_gnd_net_\,
            in3 => \N__18719\,
            lcout => \Lab_UT.dictrl.N_189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__20883\,
            in1 => \N__14800\,
            in2 => \N__14783\,
            in3 => \N__21098\,
            lcout => \Lab_UT.dictrl.state_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => \N__15871\,
            sr => \N__19207\
        );

    \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__14802\,
            in1 => \N__21021\,
            in2 => \N__14782\,
            in3 => \N__20885\,
            lcout => \Lab_UT.dictrl.state_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => \N__15871\,
            sr => \N__19207\
        );

    \Lab_UT.dictrl.state_0_esr_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__20884\,
            in1 => \N__14801\,
            in2 => \N__14784\,
            in3 => \N__21099\,
            lcout => \Lab_UT.dictrl.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => \N__15871\,
            sr => \N__19207\
        );

    \Lab_UT.dictrl.state_ret_11_RNITTE7F_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__14799\,
            in1 => \N__21020\,
            in2 => \N__14781\,
            in3 => \N__20882\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_1\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__18302\,
            in1 => \N__21097\,
            in2 => \N__14751\,
            in3 => \N__16179\,
            lcout => \Lab_UT.LdStens_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => \N__15871\,
            sr => \N__19207\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_12_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001001111"
        )
    port map (
            in0 => \N__16271\,
            in1 => \N__14853\,
            in2 => \N__14738\,
            in3 => \N__16159\,
            lcout => \Lab_UT.dictrl.N_81_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_10_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000000000"
        )
    port map (
            in0 => \N__16272\,
            in1 => \N__16283\,
            in2 => \N__14739\,
            in3 => \N__14837\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_95_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_6_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__21048\,
            in1 => \N__20906\,
            in2 => \N__14712\,
            in3 => \N__14859\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111011"
        )
    port map (
            in0 => \N__20907\,
            in1 => \N__16301\,
            in2 => \N__14709\,
            in3 => \N__16386\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__14700\,
            in1 => \N__18198\,
            in2 => \N__14706\,
            in3 => \N__14910\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000110"
        )
    port map (
            in0 => \N__18999\,
            in1 => \N__21049\,
            in2 => \N__14703\,
            in3 => \N__15583\,
            lcout => \Lab_UT.dictrl.un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18684\,
            in1 => \N__21022\,
            in2 => \N__21255\,
            in3 => \N__19802\,
            lcout => \Lab_UT.dictrl.g2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_2_5_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__16469\,
            in1 => \N__16434\,
            in2 => \N__14901\,
            in3 => \N__16781\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIQOJQ3_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__16378\,
            in1 => \N__16560\,
            in2 => \N__14880\,
            in3 => \N__18944\,
            lcout => \Lab_UT.dictrl.g2_0\,
            ltout => \Lab_UT.dictrl.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_9_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__19395\,
            in1 => \N__14868\,
            in2 => \N__14862\,
            in3 => \N__18747\,
            lcout => \Lab_UT.dictrl.N_90_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_15_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__18945\,
            in1 => \N__18786\,
            in2 => \N__16746\,
            in3 => \N__18375\,
            lcout => \Lab_UT.dictrl.m40_N_5_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__16780\,
            in1 => \N__14900\,
            in2 => \_gnd_net_\,
            in3 => \N__18943\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNI416J3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111011"
        )
    port map (
            in0 => \N__18787\,
            in1 => \N__16270\,
            in2 => \N__14847\,
            in3 => \N__16379\,
            lcout => \Lab_UT.dictrl.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIVJEO_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19376\,
            in1 => \N__20375\,
            in2 => \N__21091\,
            in3 => \N__18382\,
            lcout => \Lab_UT.dictrl.g0_17_a6_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIE4AI_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14826\,
            in1 => \N__16377\,
            in2 => \N__21092\,
            in3 => \N__18383\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFEKI3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__14820\,
            in1 => \N__14811\,
            in2 => \N__14805\,
            in3 => \N__18441\,
            lcout => \Lab_UT.dictrl.g0_17_0\,
            ltout => \Lab_UT.dictrl.g0_17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14913\,
            in3 => \N__16060\,
            lcout => \Lab_UT.dictrl.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18310\,
            in2 => \_gnd_net_\,
            in3 => \N__21057\,
            lcout => \Lab_UT.dictrl.state_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21593\,
            ce => \N__15873\,
            sr => \N__19212\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__21056\,
            in1 => \_gnd_net_\,
            in2 => \N__18315\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_dictrl_state_3_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21593\,
            ce => \N__15873\,
            sr => \N__19212\
        );

    \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18314\,
            in2 => \_gnd_net_\,
            in3 => \N__21058\,
            lcout => \Lab_UT.dictrl.state_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21593\,
            ce => \N__15873\,
            sr => \N__19212\
        );

    \buart.Z_rx.shifter_4_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20577\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21592\,
            ce => \N__19313\,
            sr => \N__19238\
        );

    \buart.Z_rx.shifter_3_rep1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20012\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21592\,
            ce => \N__19313\,
            sr => \N__19238\
        );

    \buart.Z_rx.shifter_fast_4_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20578\,
            lcout => bu_rx_data_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21592\,
            ce => \N__19313\,
            sr => \N__19238\
        );

    \buart.Z_rx.shifter_fast_3_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20013\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21592\,
            ce => \N__19313\,
            sr => \N__19238\
        );

    \Lab_UT.didp.ce_RNIDJKH1_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14924\,
            in2 => \_gnd_net_\,
            in3 => \N__15197\,
            lcout => \Lab_UT.didp.un1_dicLdMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_3_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15018\,
            in1 => \N__15959\,
            in2 => \N__15227\,
            in3 => \N__16652\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15955\,
            in1 => \N__16651\,
            in2 => \N__15226\,
            in3 => \N__15014\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15069\,
            in1 => \N__15063\,
            in2 => \N__15027\,
            in3 => \N__15477\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.ce_2_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15956\,
            in1 => \N__15219\,
            in2 => \_gnd_net_\,
            in3 => \N__15016\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.reset_1_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15017\,
            in1 => \N__15218\,
            in2 => \_gnd_net_\,
            in3 => \N__15958\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.reset_0_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15015\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.reset_2_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15019\,
            in1 => \N__15960\,
            in2 => \N__15228\,
            in3 => \N__16653\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21670\,
            ce => 'H',
            sr => \N__19214\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_3_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15430\,
            in1 => \N__15631\,
            in2 => \_gnd_net_\,
            in3 => \N__15380\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__15901\,
            in1 => \N__15341\,
            in2 => \N__14937\,
            in3 => \N__20507\,
            lcout => \Lab_UT.didp.countrce2.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100001"
        )
    port map (
            in0 => \N__14934\,
            in1 => \N__15118\,
            in2 => \N__14928\,
            in3 => \N__15198\,
            lcout => \Lab_UT.didp.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__15432\,
            in1 => \N__15340\,
            in2 => \N__15387\,
            in3 => \N__15632\,
            lcout => \Lab_UT.didp.un24_ce_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_1_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__15381\,
            in1 => \N__20298\,
            in2 => \N__15903\,
            in3 => \N__15433\,
            lcout => \Lab_UT.didp.countrce2.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__15897\,
            in1 => \N__15431\,
            in2 => \_gnd_net_\,
            in3 => \N__19928\,
            lcout => \Lab_UT.didp.countrce2.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20499\,
            in1 => \N__15189\,
            in2 => \N__15153\,
            in3 => \N__15468\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15469\,
            in1 => \N__15136\,
            in2 => \N__15105\,
            in3 => \N__15102\,
            lcout => \Lab_UT.didp.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__15379\,
            in1 => \N__15282\,
            in2 => \N__15260\,
            in3 => \N__15078\,
            lcout => \Lab_UT.didp.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16898\,
            in1 => \N__17039\,
            in2 => \_gnd_net_\,
            in3 => \N__16992\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20498\,
            in1 => \N__16942\,
            in2 => \N__15072\,
            in3 => \N__17076\,
            lcout => \Lab_UT.didp.countrce3.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15413\,
            in2 => \_gnd_net_\,
            in3 => \N__15378\,
            lcout => \Lab_UT.didp.countrce2.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI5AJE1_3_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__17337\,
            in1 => \N__17075\,
            in2 => \N__16627\,
            in3 => \N__15467\,
            lcout => \Lab_UT.didp.did_alarmMatch_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__15450\,
            in1 => \N__15252\,
            in2 => \N__15288\,
            in3 => \N__15342\,
            lcout => \Lab_UT.didp.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__15286\,
            in1 => \N__15444\,
            in2 => \N__15434\,
            in3 => \N__15259\,
            lcout => \Lab_UT.didp.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__16879\,
            in1 => \N__17452\,
            in2 => \N__16996\,
            in3 => \N__17421\,
            lcout => \Lab_UT.didp.regrce3.did_alarmMatch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__15385\,
            in1 => \N__15617\,
            in2 => \N__16815\,
            in3 => \N__17560\,
            lcout => \Lab_UT.didp.did_alarmMatch_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNITLJB1_3_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17535\,
            in1 => \N__15986\,
            in2 => \N__17263\,
            in3 => \N__15338\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.did_alarmMatch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNI08DN5_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15312\,
            in1 => \N__15306\,
            in2 => \N__15300\,
            in3 => \N__15297\,
            lcout => \Lab_UT.did_alarmMatch_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__15594\,
            in1 => \N__15287\,
            in2 => \N__15261\,
            in3 => \N__15618\,
            lcout => \Lab_UT.didp.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__17825\,
            in1 => \N__19288\,
            in2 => \_gnd_net_\,
            in3 => \N__17756\,
            lcout => \G_184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIUNGG1_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17284\,
            in1 => \N__17308\,
            in2 => \N__17956\,
            in3 => \N__16030\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.did_alarmMatch_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIO6DH5_0_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17142\,
            in1 => \N__15690\,
            in2 => \N__15678\,
            in3 => \N__15675\,
            lcout => \Lab_UT.did_alarmMatch_13\,
            ltout => \Lab_UT.did_alarmMatch_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_0__m3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__17700\,
            in1 => \N__17824\,
            in2 => \N__15669\,
            in3 => \N__15653\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__17826\,
            in2 => \N__15666\,
            in3 => \N__15493\,
            lcout => \G_183\,
            ltout => \G_183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17757\,
            in1 => \N__15663\,
            in2 => \N__15657\,
            in3 => \N__15654\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20739\,
            in1 => \N__15642\,
            in2 => \N__15902\,
            in3 => \N__15627\,
            lcout => \Lab_UT.didp.countrce2.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_armed_4_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17813\,
            in1 => \N__15578\,
            in2 => \_gnd_net_\,
            in3 => \N__17736\,
            lcout => \Lab_UT.alarmstate_0_sqmuxa_1\,
            ltout => \Lab_UT.alarmstate_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_idle_5_0_iclk_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110001"
        )
    port map (
            in0 => \N__17738\,
            in1 => \N__17815\,
            in2 => \N__15516\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.un1_idle_5_0_iclkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__17755\,
            in1 => \N__15513\,
            in2 => \N__15501\,
            in3 => \N__17640\,
            lcout => \G_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__15852\,
            in1 => \N__20740\,
            in2 => \N__18002\,
            in3 => \N__16043\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__15801\,
            in1 => \N__16039\,
            in2 => \N__15846\,
            in3 => \N__15832\,
            lcout => \Lab_UT.didp.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__15831\,
            in1 => \N__17910\,
            in2 => \N__17960\,
            in3 => \N__15802\,
            lcout => \Lab_UT.didp.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.un1_armed_2_0_iso_i_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17737\,
            lcout => \Lab_UT.un1_armed_2_0_iso_iZ0\,
            ltout => \Lab_UT.un1_armed_2_0_iso_iZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_latch_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__15765\,
            in1 => \N__15751\,
            in2 => \N__15708\,
            in3 => \N__15705\,
            lcout => \G_192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__21103\,
            in1 => \N__18186\,
            in2 => \_gnd_net_\,
            in3 => \N__17859\,
            lcout => \Lab_UT.dictrl.state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => \N__15869\,
            sr => \N__19205\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19527\,
            in1 => \N__17877\,
            in2 => \_gnd_net_\,
            in3 => \N__19756\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__21101\,
            in2 => \N__15693\,
            in3 => \N__20893\,
            lcout => \Lab_UT.state_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => \N__15869\,
            sr => \N__19205\
        );

    \Lab_UT.dictrl.state_0_esr_2_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17896\,
            in1 => \N__16115\,
            in2 => \N__18177\,
            in3 => \N__16082\,
            lcout => \Lab_UT.dictrl.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => \N__15869\,
            sr => \N__19205\
        );

    \Lab_UT.dictrl.state_0_fast_esr_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__16083\,
            in1 => \N__18174\,
            in2 => \N__16119\,
            in3 => \N__17897\,
            lcout => \Lab_UT.dictrl.state_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => \N__15869\,
            sr => \N__19205\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17895\,
            in1 => \N__16114\,
            in2 => \N__18176\,
            in3 => \N__16081\,
            lcout => \Lab_UT.dictrl.state_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => \N__15869\,
            sr => \N__19205\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNIAD6S_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21197\,
            in1 => \N__18253\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => \Lab_UT.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16034\,
            in1 => \N__17949\,
            in2 => \N__18068\,
            in3 => \N__15998\,
            lcout => \Lab_UT.didp.un18_ce\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__16177\,
            in1 => \N__18297\,
            in2 => \_gnd_net_\,
            in3 => \N__21083\,
            lcout => \Lab_UT.LdSones_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21621\,
            ce => \N__15870\,
            sr => \N__19208\
        );

    \Lab_UT.dictrl.state_ret_4_esr_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21079\,
            in1 => \N__18287\,
            in2 => \_gnd_net_\,
            in3 => \N__16176\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21621\,
            ce => \N__15870\,
            sr => \N__19208\
        );

    \Lab_UT.dictrl.state_0_esr_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16188\,
            in1 => \N__18542\,
            in2 => \N__21102\,
            in3 => \N__20887\,
            lcout => \Lab_UT.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21621\,
            ce => \N__15870\,
            sr => \N__19208\
        );

    \Lab_UT.dictrl.state_ret_6_esr_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__16178\,
            in1 => \N__15917\,
            in2 => \N__18298\,
            in3 => \N__21084\,
            lcout => \Lab_UT.LdStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21621\,
            ce => \N__15870\,
            sr => \N__19208\
        );

    \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21078\,
            in2 => \_gnd_net_\,
            in3 => \N__18286\,
            lcout => \Lab_UT.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21621\,
            ce => \N__15870\,
            sr => \N__19208\
        );

    \Lab_UT.dictrl.m25_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__16534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18912\,
            lcout => \Lab_UT.dictrl.m25Z0Z_0\,
            ltout => \Lab_UT.dictrl.m25Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m30_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16407\,
            in1 => \N__16227\,
            in2 => \N__16206\,
            in3 => \N__20380\,
            lcout => \Lab_UT.dictrl.N_114_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m59_ns_1_x1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__16533\,
            in1 => \N__18911\,
            in2 => \N__18605\,
            in3 => \N__16406\,
            lcout => \Lab_UT.dictrl.m59_ns_1_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_RNILO8G6_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100000101"
        )
    port map (
            in0 => \N__16160\,
            in1 => \N__19420\,
            in2 => \N__18750\,
            in3 => \N__17586\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_81_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIB544A_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19520\,
            in2 => \N__16191\,
            in3 => \N__19794\,
            lcout => \Lab_UT.dictrl.N_113_1\,
            ltout => \Lab_UT.dictrl.N_113_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNIC32CN_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20881\,
            in1 => \N__21023\,
            in2 => \N__16182\,
            in3 => \N__18543\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNITSVD3_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__19421\,
            in1 => \N__18104\,
            in2 => \_gnd_net_\,
            in3 => \N__19793\,
            lcout => \Lab_UT.dictrl.i10_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNII0R67_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110101"
        )
    port map (
            in0 => \N__19645\,
            in1 => \N__21196\,
            in2 => \N__18108\,
            in3 => \N__16161\,
            lcout => \Lab_UT.dictrl.N_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m40_m2_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__18789\,
            in1 => \N__21324\,
            in2 => \N__20254\,
            in3 => \N__18846\,
            lcout => \Lab_UT.dictrl.m40_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m73_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21325\,
            in1 => \N__20753\,
            in2 => \_gnd_net_\,
            in3 => \N__19912\,
            lcout => \Lab_UT.dictrl.m73Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_11_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19407\,
            in2 => \_gnd_net_\,
            in3 => \N__18749\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_16_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_7_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__19795\,
            in1 => \N__16395\,
            in2 => \N__16389\,
            in3 => \N__16662\,
            lcout => \Lab_UT.dictrl.N_113_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_23_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__16233\,
            in1 => \N__18850\,
            in2 => \N__16751\,
            in3 => \N__18354\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNI1N6L5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111100000110"
        )
    port map (
            in0 => \N__18748\,
            in1 => \N__16366\,
            in2 => \N__16317\,
            in3 => \N__16551\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNI5EFJC_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__16314\,
            in1 => \N__16542\,
            in2 => \N__16308\,
            in3 => \N__19408\,
            lcout => \Lab_UT.dictrl.i9_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_12_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__18353\,
            in1 => \N__18788\,
            in2 => \N__18866\,
            in3 => \N__16745\,
            lcout => \Lab_UT.dictrl.N_77_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_16_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100101111"
        )
    port map (
            in0 => \N__16260\,
            in1 => \N__18851\,
            in2 => \N__16752\,
            in3 => \N__18355\,
            lcout => \Lab_UT.dictrl.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__16433\,
            in1 => \N__16531\,
            in2 => \N__16485\,
            in3 => \N__18901\,
            lcout => \Lab_UT.dictrl.g0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_2_4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__18900\,
            in1 => \_gnd_net_\,
            in2 => \N__16536\,
            in3 => \N__18419\,
            lcout => \Lab_UT.dictrl.g0_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_4_2_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__16484\,
            in1 => \N__18940\,
            in2 => \N__16785\,
            in3 => \N__16532\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_22_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19498\,
            in1 => \N__16750\,
            in2 => \N__16554\,
            in3 => \N__20573\,
            lcout => \Lab_UT.dictrl.N_77_1_0\,
            ltout => \Lab_UT.dictrl.N_77_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNI11N26_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__19396\,
            in1 => \N__16680\,
            in2 => \N__16545\,
            in3 => \N__18515\,
            lcout => \Lab_UT.dictrl.N_2353_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m37_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18899\,
            in1 => \N__16479\,
            in2 => \N__16535\,
            in3 => \N__16432\,
            lcout => \Lab_UT.dictrl.N_103_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIQTDF1_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__16480\,
            in1 => \N__16455\,
            in2 => \N__18910\,
            in3 => \N__16779\,
            lcout => \Lab_UT.dictrl.g1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m47_x0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16423\,
            in1 => \N__20157\,
            in2 => \N__18628\,
            in3 => \N__20570\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m47_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m47_ns_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16437\,
            in3 => \N__16778\,
            lcout => \Lab_UT.dictrl.N_106_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m30_1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16422\,
            in2 => \_gnd_net_\,
            in3 => \N__16777\,
            lcout => \Lab_UT.dictrl.m30Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_1_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20754\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__19314\,
            sr => \N__19239\
        );

    \buart.Z_rx.shifter_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20158\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__19314\,
            sr => \N__19239\
        );

    \Lab_UT.dictrl.g1_1_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16720\,
            in1 => \N__18423\,
            in2 => \_gnd_net_\,
            in3 => \N__18874\,
            lcout => \Lab_UT.dictrl.g1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__20003\,
            in1 => \N__16671\,
            in2 => \_gnd_net_\,
            in3 => \N__18570\,
            lcout => \Lab_UT.dictrl.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17049\,
            in1 => \N__17002\,
            in2 => \N__16905\,
            in3 => \N__17087\,
            lcout => \Lab_UT.didp.countrce3.ce_12_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_0_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19956\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21671\,
            ce => \N__16605\,
            sr => \N__19215\
        );

    \Lab_UT.didp.regrce4.q_esr_3_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20508\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21671\,
            ce => \N__16605\,
            sr => \N__19215\
        );

    \Lab_UT.didp.ce_RNI4EIS1_2_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17231\,
            in2 => \_gnd_net_\,
            in3 => \N__16955\,
            lcout => \Lab_UT.didp.un1_dicLdMones_0\,
            ltout => \Lab_UT.didp.un1_dicLdMones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__16991\,
            in1 => \N__17127\,
            in2 => \N__16575\,
            in3 => \N__16572\,
            lcout => \Lab_UT.didp.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001001"
        )
    port map (
            in0 => \N__17232\,
            in1 => \N__17217\,
            in2 => \N__17130\,
            in3 => \N__16956\,
            lcout => \Lab_UT.didp.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__16900\,
            in1 => \N__17128\,
            in2 => \N__16857\,
            in3 => \N__17096\,
            lcout => \Lab_UT.didp.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__17027\,
            in1 => \N__17197\,
            in2 => \N__17503\,
            in3 => \N__17158\,
            lcout => \Lab_UT.didp.regrce4.did_alarmMatch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17083\,
            in1 => \N__17129\,
            in2 => \N__17106\,
            in3 => \N__17097\,
            lcout => \Lab_UT.didp.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16990\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__16954\,
            in1 => \N__20741\,
            in2 => \N__16908\,
            in3 => \N__16899\,
            lcout => \Lab_UT.didp.countrce3.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__20925\,
            in1 => \N__16842\,
            in2 => \N__17400\,
            in3 => \N__19950\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce2.q_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__20926\,
            in2 => \N__16822\,
            in3 => \N__17387\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce2.q_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__20927\,
            in1 => \N__20742\,
            in2 => \N__17401\,
            in3 => \N__17566\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce2.q_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20496\,
            in1 => \N__20928\,
            in2 => \N__17542\,
            in3 => \N__17391\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce3.q_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__17630\,
            in1 => \N__17493\,
            in2 => \N__17402\,
            in3 => \N__19951\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce3.q_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20297\,
            in1 => \N__17631\,
            in2 => \N__17464\,
            in3 => \N__17395\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce3.q_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__17632\,
            in1 => \N__20743\,
            in2 => \N__17403\,
            in3 => \N__17428\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce3.q_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20497\,
            in1 => \N__17633\,
            in2 => \N__17353\,
            in3 => \N__17399\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21658\,
            ce => 'H',
            sr => \N__19213\
        );

    \Lab_UT.didp.regrce1.q_esr_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20295\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21652\,
            ce => \N__18662\,
            sr => \N__19211\
        );

    \Lab_UT.didp.regrce1.q_esr_2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20731\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21652\,
            ce => \N__18662\,
            sr => \N__19211\
        );

    \Lab_UT.didp.regrce1.q_esr_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20492\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21652\,
            ce => \N__18662\,
            sr => \N__19211\
        );

    \Lab_UT.dictrl.alarmstate8_3_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19499\,
            in1 => \N__20168\,
            in2 => \N__20609\,
            in3 => \N__19905\,
            lcout => \Lab_UT.dictrl.alarmstate8Z0Z_3\,
            ltout => \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_0__m3_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__17827\,
            in1 => \N__17767\,
            in2 => \N__17703\,
            in3 => \N__18077\,
            lcout => \Lab_UT.dictrl.m3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.justentered_1_sqmuxa_i_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__17651\,
            in1 => \N__17676\,
            in2 => \N__17670\,
            in3 => \N__19289\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.justentered_latch_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__17691\,
            in1 => \_gnd_net_\,
            in2 => \N__17694\,
            in3 => \N__17652\,
            lcout => \G_188\,
            ltout => \G_188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate22_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__17685\,
            in1 => \_gnd_net_\,
            in2 => \N__17679\,
            in3 => \N__18078\,
            lcout => \G_187\,
            ltout => \G_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17669\,
            in2 => \N__17655\,
            in3 => \N__17650\,
            lcout => \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIA8O21_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21251\,
            in1 => \N__18493\,
            in2 => \N__17629\,
            in3 => \N__19739\,
            lcout => \Lab_UT.LdASones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_2_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__19503\,
            in1 => \N__20156\,
            in2 => \N__18632\,
            in3 => \N__20602\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_15_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__18854\,
            in1 => \N__18379\,
            in2 => \N__17589\,
            in3 => \N__21333\,
            lcout => \Lab_UT.dictrl.m40_N_5_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate8_4_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18853\,
            in1 => \N__20379\,
            in2 => \N__18384\,
            in3 => \N__21332\,
            lcout => \Lab_UT.dictrl.alarmstate8Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20285\,
            in1 => \N__18069\,
            in2 => \N__17994\,
            in3 => \N__17952\,
            lcout => \Lab_UT.didp.countrce1.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21628\,
            ce => \N__19319\,
            sr => \N__19236\
        );

    \Lab_UT.dictrl.g0_17_o3_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20427\,
            in2 => \_gnd_net_\,
            in3 => \N__20671\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIS3A93_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110101"
        )
    port map (
            in0 => \N__20879\,
            in1 => \N__18798\,
            in2 => \N__17904\,
            in3 => \N__19676\,
            lcout => \Lab_UT.dictrl.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20426\,
            in2 => \_gnd_net_\,
            in3 => \N__20670\,
            lcout => \Lab_UT.dictrl.m51_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__20880\,
            in1 => \N__18450\,
            in2 => \N__17876\,
            in3 => \N__19755\,
            lcout => \Lab_UT.dictrl.next_state_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20057\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21628\,
            ce => \N__19319\,
            sr => \N__19236\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_5_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110101010101"
        )
    port map (
            in0 => \N__19655\,
            in1 => \N__18264\,
            in2 => \N__18144\,
            in3 => \N__20038\,
            lcout => \Lab_UT.dictrl.P8_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUI6O8_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__20878\,
            in1 => \N__18219\,
            in2 => \N__18213\,
            in3 => \N__18135\,
            lcout => \Lab_UT.dictrl.next_state_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_12_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110111"
        )
    port map (
            in0 => \N__20264\,
            in1 => \N__20698\,
            in2 => \N__19809\,
            in3 => \N__20472\,
            lcout => \Lab_UT.dictrl.P6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNI0C4D4_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__18257\,
            in1 => \N__19419\,
            in2 => \N__18231\,
            in3 => \N__19654\,
            lcout => \Lab_UT.dictrl.N_69\,
            ltout => \Lab_UT.dictrl.N_69_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__18134\,
            in1 => \N__18212\,
            in2 => \N__18201\,
            in3 => \N__20877\,
            lcout => \Lab_UT.dictrl.next_state_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19781\,
            in1 => \N__18090\,
            in2 => \N__19677\,
            in3 => \N__20775\,
            lcout => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNIIOLT_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__21176\,
            in2 => \_gnd_net_\,
            in3 => \N__19780\,
            lcout => \Lab_UT.dictrl.g0_17_a6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_11_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101110101"
        )
    port map (
            in0 => \N__20471\,
            in1 => \N__20697\,
            in2 => \N__21216\,
            in3 => \N__20263\,
            lcout => \Lab_UT.dictrl.P6_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI00K56_3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__18133\,
            in1 => \N__18089\,
            in2 => \N__21238\,
            in3 => \N__18103\,
            lcout => \Lab_UT.dictrl.m77_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m55_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__20250\,
            in1 => \N__18790\,
            in2 => \N__20764\,
            in3 => \N__21326\,
            lcout => \Lab_UT.dictrl.N_77\,
            ltout => \Lab_UT.dictrl.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIRLAN5_3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__18522\,
            in1 => \N__21211\,
            in2 => \N__18564\,
            in3 => \N__18561\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIASHNC_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__18552\,
            in1 => \N__19672\,
            in2 => \N__18546\,
            in3 => \N__19778\,
            lcout => \Lab_UT.dictrl.i9_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__18521\,
            in1 => \N__18504\,
            in2 => \N__21239\,
            in3 => \N__19927\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_118_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111000000"
        )
    port map (
            in0 => \N__21212\,
            in1 => \N__18495\,
            in2 => \N__18453\,
            in3 => \N__19779\,
            lcout => \Lab_UT.dictrl.next_state_latmux_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_17_a6_3_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20155\,
            in1 => \N__20604\,
            in2 => \N__20052\,
            in3 => \N__19926\,
            lcout => \Lab_UT.dictrl.g0_17_a6_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_fast_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20246\,
            lcout => \buart__rx_shifter_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_1_rep1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_2_rep1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20488\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_fast_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_3_rep2_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20048\,
            lcout => bu_rx_data_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \buart.Z_rx.shifter_fast_5_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20160\,
            lcout => \buart__rx_shifter_fast_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => \N__19317\,
            sr => \N__19240\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_RNID53P_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19402\,
            in2 => \_gnd_net_\,
            in3 => \N__18751\,
            lcout => \N_16_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_8_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18852\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_11_RNO_5_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110101"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__18791\,
            in2 => \N__18756\,
            in3 => \N__18752\,
            lcout => \Lab_UT.dictrl.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_rep2_RNIT8A31_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011011111"
        )
    port map (
            in0 => \N__20223\,
            in1 => \N__19403\,
            in2 => \N__20755\,
            in3 => \N__21327\,
            lcout => \buart.Z_rx.P7_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18672\,
            in2 => \_gnd_net_\,
            in3 => \N__19285\,
            lcout => \Lab_UT.didp.regrce1.LdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_rep1_RNIG7Q01_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18627\,
            in1 => \N__20159\,
            in2 => \_gnd_net_\,
            in3 => \N__20571\,
            lcout => \shifter_7_rep1_RNIG7Q01\,
            ltout => \shifter_7_rep1_RNIG7Q01_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIUOH63_4_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__19536\,
            in2 => \N__19530\,
            in3 => \N__20030\,
            lcout => \N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_rep1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20572\,
            lcout => bu_rx_data_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21597\,
            ce => \N__19315\,
            sr => \N__19241\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_ctle_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19017\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19283\,
            lcout => bu_rx_data_rdy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_9_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19812\,
            in1 => \N__20169\,
            in2 => \N__19428\,
            in3 => \N__19873\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_5_a4_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__21276\,
            in1 => \N__20056\,
            in2 => \N__19338\,
            in3 => \N__20287\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__21236\,
            in1 => \N__19554\,
            in2 => \N__19335\,
            in3 => \N__19671\,
            lcout => \Lab_UT.dictrl.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21639\,
            ce => \N__19320\,
            sr => \N__19237\
        );

    \Lab_UT.dictrl.m86_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19010\,
            in1 => \N__21267\,
            in2 => \N__18960\,
            in3 => \N__20388\,
            lcout => \N_119_mux\,
            ltout => \N_119_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21398\,
            in2 => \N__21360\,
            in3 => \N__21759\,
            lcout => \resetGen_reset_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_8_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20610\,
            in1 => \N__20757\,
            in2 => \N__21357\,
            in3 => \N__20387\,
            lcout => \Lab_UT.dictrl.g0_5_a4_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m86_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20037\,
            in2 => \_gnd_net_\,
            in3 => \N__20284\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m86Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m86_2_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20490\,
            in1 => \N__20756\,
            in2 => \N__21270\,
            in3 => \N__19872\,
            lcout => \Lab_UT.dictrl.m86Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21243\,
            in1 => \N__21105\,
            in2 => \_gnd_net_\,
            in3 => \N__20936\,
            lcout => \Lab_UT.dictrl.next_state_latmux_1_a0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_6_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__20603\,
            in2 => \N__20506\,
            in3 => \N__20373\,
            lcout => \Lab_UT.dictrl.g0_5_o4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_7_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__20286\,
            in1 => \N__20162\,
            in2 => \N__20058\,
            in3 => \N__19888\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_5_o4_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__19821\,
            in1 => \N__19811\,
            in2 => \N__19680\,
            in3 => \N__19670\,
            lcout => \Lab_UT.dictrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m90_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21417\,
            in1 => \N__21755\,
            in2 => \N__21713\,
            in3 => \N__21729\,
            lcout => \N_91_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m93_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__21757\,
            in1 => \N__21419\,
            in2 => \N__21737\,
            in3 => \N__21711\,
            lcout => OPEN,
            ltout => \N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__21689\,
            in1 => \N__21366\,
            in2 => \N__21762\,
            in3 => \N__21680\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010010"
        )
    port map (
            in0 => \N__21758\,
            in1 => \N__21421\,
            in2 => \N__21738\,
            in3 => \N__21392\,
            lcout => \resetGen_reset_count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m97_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__21418\,
            in1 => \N__21756\,
            in2 => \N__21714\,
            in3 => \N__21730\,
            lcout => OPEN,
            ltout => \resetGen_reset_count_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__21396\,
            in1 => \N__21423\,
            in2 => \N__21717\,
            in3 => \N__21712\,
            lcout => \resetGen_reset_count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__21422\,
            in1 => \N__21397\,
            in2 => \N__21693\,
            in3 => \N__21681\,
            lcout => \resetGen_reset_count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m87_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21420\,
            in2 => \_gnd_net_\,
            in3 => \N__21391\,
            lcout => m87,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
